magic
tech sky130A
magscale 1 2
timestamp 1654688367
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 314654 700952 314660 701004
rect 314712 700992 314718 701004
rect 413646 700992 413652 701004
rect 314712 700964 413652 700992
rect 314712 700952 314718 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 325694 700884 325700 700936
rect 325752 700924 325758 700936
rect 429838 700924 429844 700936
rect 325752 700896 429844 700924
rect 325752 700884 325758 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 336734 700816 336740 700868
rect 336792 700856 336798 700868
rect 446122 700856 446128 700868
rect 336792 700828 446128 700856
rect 336792 700816 336798 700828
rect 446122 700816 446128 700828
rect 446180 700816 446186 700868
rect 347866 700748 347872 700800
rect 347924 700788 347930 700800
rect 462314 700788 462320 700800
rect 347924 700760 462320 700788
rect 347924 700748 347930 700760
rect 462314 700748 462320 700760
rect 462372 700748 462378 700800
rect 358814 700680 358820 700732
rect 358872 700720 358878 700732
rect 478506 700720 478512 700732
rect 358872 700692 478512 700720
rect 358872 700680 358878 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 248414 700612 248420 700664
rect 248472 700652 248478 700664
rect 316310 700652 316316 700664
rect 248472 700624 316316 700652
rect 248472 700612 248478 700624
rect 316310 700612 316316 700624
rect 316368 700612 316374 700664
rect 369854 700612 369860 700664
rect 369912 700652 369918 700664
rect 494790 700652 494796 700664
rect 369912 700624 494796 700652
rect 369912 700612 369918 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 259454 700544 259460 700596
rect 259512 700584 259518 700596
rect 332502 700584 332508 700596
rect 259512 700556 332508 700584
rect 259512 700544 259518 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 379514 700544 379520 700596
rect 379572 700584 379578 700596
rect 510982 700584 510988 700596
rect 379572 700556 510988 700584
rect 379572 700544 379578 700556
rect 510982 700544 510988 700556
rect 511040 700544 511046 700596
rect 204254 700476 204260 700528
rect 204312 700516 204318 700528
rect 251450 700516 251456 700528
rect 204312 700488 251456 700516
rect 204312 700476 204318 700488
rect 251450 700476 251456 700488
rect 251508 700476 251514 700528
rect 270494 700476 270500 700528
rect 270552 700516 270558 700528
rect 348786 700516 348792 700528
rect 270552 700488 348792 700516
rect 270552 700476 270558 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 390554 700476 390560 700528
rect 390612 700516 390618 700528
rect 527174 700516 527180 700528
rect 390612 700488 527180 700516
rect 390612 700476 390618 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 171134 700408 171140 700460
rect 171192 700448 171198 700460
rect 202782 700448 202788 700460
rect 171192 700420 202788 700448
rect 171192 700408 171198 700420
rect 202782 700408 202788 700420
rect 202840 700408 202846 700460
rect 215294 700408 215300 700460
rect 215352 700448 215358 700460
rect 267642 700448 267648 700460
rect 215352 700420 267648 700448
rect 215352 700408 215358 700420
rect 267642 700408 267648 700420
rect 267700 700408 267706 700460
rect 281534 700408 281540 700460
rect 281592 700448 281598 700460
rect 364978 700448 364984 700460
rect 281592 700420 364984 700448
rect 281592 700408 281598 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 401594 700408 401600 700460
rect 401652 700448 401658 700460
rect 543458 700448 543464 700460
rect 401652 700420 543464 700448
rect 401652 700408 401658 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 149054 700340 149060 700392
rect 149112 700380 149118 700392
rect 170306 700380 170312 700392
rect 149112 700352 170312 700380
rect 149112 700340 149118 700352
rect 170306 700340 170312 700352
rect 170364 700340 170370 700392
rect 182174 700340 182180 700392
rect 182232 700380 182238 700392
rect 218974 700380 218980 700392
rect 182232 700352 218980 700380
rect 182232 700340 182238 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 226334 700340 226340 700392
rect 226392 700380 226398 700392
rect 283834 700380 283840 700392
rect 226392 700352 283840 700380
rect 226392 700340 226398 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 292574 700340 292580 700392
rect 292632 700380 292638 700392
rect 381170 700380 381176 700392
rect 292632 700352 381176 700380
rect 292632 700340 292638 700352
rect 381170 700340 381176 700352
rect 381228 700340 381234 700392
rect 412634 700340 412640 700392
rect 412692 700380 412698 700392
rect 559650 700380 559656 700392
rect 412692 700352 559656 700380
rect 412692 700340 412698 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 126974 700272 126980 700324
rect 127032 700312 127038 700324
rect 137830 700312 137836 700324
rect 127032 700284 137836 700312
rect 127032 700272 127038 700284
rect 137830 700272 137836 700284
rect 137888 700272 137894 700324
rect 138014 700272 138020 700324
rect 138072 700312 138078 700324
rect 154114 700312 154120 700324
rect 138072 700284 154120 700312
rect 138072 700272 138078 700284
rect 154114 700272 154120 700284
rect 154172 700272 154178 700324
rect 160094 700272 160100 700324
rect 160152 700312 160158 700324
rect 186498 700312 186504 700324
rect 160152 700284 186504 700312
rect 160152 700272 160158 700284
rect 186498 700272 186504 700284
rect 186556 700272 186562 700324
rect 193214 700272 193220 700324
rect 193272 700312 193278 700324
rect 235166 700312 235172 700324
rect 193272 700284 235172 700312
rect 193272 700272 193278 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 237374 700272 237380 700324
rect 237432 700312 237438 700324
rect 300118 700312 300124 700324
rect 237432 700284 300124 700312
rect 237432 700272 237438 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 303614 700272 303620 700324
rect 303672 700312 303678 700324
rect 397454 700312 397460 700324
rect 303672 700284 397460 700312
rect 303672 700272 303678 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 423674 700272 423680 700324
rect 423732 700312 423738 700324
rect 575842 700312 575848 700324
rect 423732 700284 575848 700312
rect 423732 700272 423738 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 115934 699660 115940 699712
rect 115992 699700 115998 699712
rect 121638 699700 121644 699712
rect 115992 699672 121644 699700
rect 115992 699660 115998 699672
rect 121638 699660 121644 699672
rect 121696 699660 121702 699712
rect 3418 683748 3424 683800
rect 3476 683788 3482 683800
rect 11698 683788 11704 683800
rect 3476 683760 11704 683788
rect 3476 683748 3482 683760
rect 11698 683748 11704 683760
rect 11756 683748 11762 683800
rect 428458 683136 428464 683188
rect 428516 683176 428522 683188
rect 579614 683176 579620 683188
rect 428516 683148 579620 683176
rect 428516 683136 428522 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3510 670964 3516 671016
rect 3568 671004 3574 671016
rect 4798 671004 4804 671016
rect 3568 670976 4804 671004
rect 3568 670964 3574 670976
rect 4798 670964 4804 670976
rect 4856 670964 4862 671016
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 33778 656928 33784 656940
rect 3568 656900 33784 656928
rect 3568 656888 3574 656900
rect 33778 656888 33784 656900
rect 33836 656888 33842 656940
rect 2866 644444 2872 644496
rect 2924 644484 2930 644496
rect 10318 644484 10324 644496
rect 2924 644456 10324 644484
rect 2924 644444 2930 644456
rect 10318 644444 10324 644456
rect 10376 644444 10382 644496
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 22738 632108 22744 632120
rect 3568 632080 22744 632108
rect 3568 632068 3574 632080
rect 22738 632068 22744 632080
rect 22796 632068 22802 632120
rect 428550 630640 428556 630692
rect 428608 630680 428614 630692
rect 579614 630680 579620 630692
rect 428608 630652 579620 630680
rect 428608 630640 428614 630652
rect 579614 630640 579620 630652
rect 579672 630640 579678 630692
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 36538 605860 36544 605872
rect 3384 605832 36544 605860
rect 3384 605820 3390 605832
rect 36538 605820 36544 605832
rect 36596 605820 36602 605872
rect 3326 592016 3332 592068
rect 3384 592056 3390 592068
rect 14458 592056 14464 592068
rect 3384 592028 14464 592056
rect 3384 592016 3390 592028
rect 14458 592016 14464 592028
rect 14516 592016 14522 592068
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 25498 579680 25504 579692
rect 3384 579652 25504 579680
rect 3384 579640 3390 579652
rect 25498 579640 25504 579652
rect 25556 579640 25562 579692
rect 428642 576852 428648 576904
rect 428700 576892 428706 576904
rect 580166 576892 580172 576904
rect 428700 576864 580172 576892
rect 428700 576852 428706 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 88334 562980 88340 563032
rect 88392 563020 88398 563032
rect 94590 563020 94596 563032
rect 88392 562992 94596 563020
rect 88392 562980 88398 562992
rect 94590 562980 94596 562992
rect 94648 562980 94654 563032
rect 40034 562436 40040 562488
rect 40092 562476 40098 562488
rect 61654 562476 61660 562488
rect 40092 562448 61660 562476
rect 40092 562436 40098 562448
rect 61654 562436 61660 562448
rect 61712 562436 61718 562488
rect 71774 562436 71780 562488
rect 71832 562476 71838 562488
rect 83642 562476 83648 562488
rect 71832 562448 83648 562476
rect 71832 562436 71838 562448
rect 83642 562436 83648 562448
rect 83700 562436 83706 562488
rect 23474 562368 23480 562420
rect 23532 562408 23538 562420
rect 50614 562408 50620 562420
rect 23532 562380 50620 562408
rect 23532 562368 23538 562380
rect 50614 562368 50620 562380
rect 50672 562368 50678 562420
rect 6914 562300 6920 562352
rect 6972 562340 6978 562352
rect 40402 562340 40408 562352
rect 6972 562312 40408 562340
rect 6972 562300 6978 562312
rect 40402 562300 40408 562312
rect 40460 562300 40466 562352
rect 56594 562300 56600 562352
rect 56652 562340 56658 562352
rect 72694 562340 72700 562352
rect 56652 562312 72700 562340
rect 56652 562300 56658 562312
rect 72694 562300 72700 562312
rect 72752 562300 72758 562352
rect 3142 553528 3148 553580
rect 3200 553568 3206 553580
rect 6178 553568 6184 553580
rect 3200 553540 6184 553568
rect 3200 553528 3206 553540
rect 6178 553528 6184 553540
rect 6236 553528 6242 553580
rect 490558 550604 490564 550656
rect 490616 550644 490622 550656
rect 580166 550644 580172 550656
rect 490616 550616 580172 550644
rect 490616 550604 490622 550616
rect 580166 550604 580172 550616
rect 580224 550604 580230 550656
rect 11698 545028 11704 545080
rect 11756 545068 11762 545080
rect 37826 545068 37832 545080
rect 11756 545040 37832 545068
rect 11756 545028 11762 545040
rect 37826 545028 37832 545040
rect 37884 545028 37890 545080
rect 428734 545028 428740 545080
rect 428792 545068 428798 545080
rect 580258 545068 580264 545080
rect 428792 545040 580264 545068
rect 428792 545028 428798 545040
rect 580258 545028 580264 545040
rect 580316 545028 580322 545080
rect 22738 541628 22744 541680
rect 22796 541668 22802 541680
rect 37918 541668 37924 541680
rect 22796 541640 37924 541668
rect 22796 541628 22802 541640
rect 37918 541628 37924 541640
rect 37976 541628 37982 541680
rect 3050 539588 3056 539640
rect 3108 539628 3114 539640
rect 22738 539628 22744 539640
rect 3108 539600 22744 539628
rect 3108 539588 3114 539600
rect 22738 539588 22744 539600
rect 22796 539588 22802 539640
rect 4798 536732 4804 536784
rect 4856 536772 4862 536784
rect 37550 536772 37556 536784
rect 4856 536744 37556 536772
rect 4856 536732 4862 536744
rect 37550 536732 37556 536744
rect 37608 536732 37614 536784
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 28258 527184 28264 527196
rect 3016 527156 28264 527184
rect 3016 527144 3022 527156
rect 28258 527144 28264 527156
rect 28316 527144 28322 527196
rect 3418 527076 3424 527128
rect 3476 527116 3482 527128
rect 37826 527116 37832 527128
rect 3476 527088 37832 527116
rect 3476 527076 3482 527088
rect 37826 527076 37832 527088
rect 37884 527076 37890 527128
rect 428734 525716 428740 525768
rect 428792 525756 428798 525768
rect 580350 525756 580356 525768
rect 428792 525728 580356 525756
rect 428792 525716 428798 525728
rect 580350 525716 580356 525728
rect 580408 525716 580414 525768
rect 428458 524424 428464 524476
rect 428516 524464 428522 524476
rect 580166 524464 580172 524476
rect 428516 524436 580172 524464
rect 428516 524424 428522 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 33778 517420 33784 517472
rect 33836 517460 33842 517472
rect 38010 517460 38016 517472
rect 33836 517432 38016 517460
rect 33836 517420 33842 517432
rect 38010 517420 38016 517432
rect 38068 517420 38074 517472
rect 428734 516060 428740 516112
rect 428792 516100 428798 516112
rect 580442 516100 580448 516112
rect 428792 516072 580448 516100
rect 428792 516060 428798 516072
rect 580442 516060 580448 516072
rect 580500 516060 580506 516112
rect 10318 507764 10324 507816
rect 10376 507804 10382 507816
rect 37550 507804 37556 507816
rect 10376 507776 37556 507804
rect 10376 507764 10382 507776
rect 37550 507764 37556 507776
rect 37608 507764 37614 507816
rect 428734 506404 428740 506456
rect 428792 506444 428798 506456
rect 580534 506444 580540 506456
rect 428792 506416 580540 506444
rect 428792 506404 428798 506416
rect 580534 506404 580540 506416
rect 580592 506404 580598 506456
rect 3142 488520 3148 488572
rect 3200 488560 3206 488572
rect 10318 488560 10324 488572
rect 3200 488532 10324 488560
rect 3200 488520 3206 488532
rect 10318 488520 10324 488532
rect 10376 488520 10382 488572
rect 3510 488452 3516 488504
rect 3568 488492 3574 488504
rect 37826 488492 37832 488504
rect 3568 488464 37832 488492
rect 3568 488452 3574 488464
rect 37826 488452 37832 488464
rect 37884 488452 37890 488504
rect 428550 487092 428556 487144
rect 428608 487132 428614 487144
rect 580626 487132 580632 487144
rect 428608 487104 580632 487132
rect 428608 487092 428614 487104
rect 580626 487092 580632 487104
rect 580684 487092 580690 487144
rect 428550 477436 428556 477488
rect 428608 477476 428614 477488
rect 580718 477476 580724 477488
rect 428608 477448 580724 477476
rect 428608 477436 428614 477448
rect 580718 477436 580724 477448
rect 580776 477436 580782 477488
rect 3510 474716 3516 474768
rect 3568 474756 3574 474768
rect 31018 474756 31024 474768
rect 3568 474728 31024 474756
rect 3568 474716 3574 474728
rect 31018 474716 31024 474728
rect 31076 474716 31082 474768
rect 428550 470568 428556 470620
rect 428608 470608 428614 470620
rect 579982 470608 579988 470620
rect 428608 470580 579988 470608
rect 428608 470568 428614 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 14458 469140 14464 469192
rect 14516 469180 14522 469192
rect 37918 469180 37924 469192
rect 14516 469152 37924 469180
rect 14516 469140 14522 469152
rect 37918 469140 37924 469152
rect 37976 469140 37982 469192
rect 428734 467780 428740 467832
rect 428792 467820 428798 467832
rect 580718 467820 580724 467832
rect 428792 467792 580724 467820
rect 428792 467780 428798 467792
rect 580718 467780 580724 467792
rect 580776 467780 580782 467832
rect 25498 459484 25504 459536
rect 25556 459524 25562 459536
rect 37458 459524 37464 459536
rect 25556 459496 37464 459524
rect 25556 459484 25562 459496
rect 37458 459484 37464 459496
rect 37516 459484 37522 459536
rect 3602 449828 3608 449880
rect 3660 449868 3666 449880
rect 37918 449868 37924 449880
rect 3660 449840 37924 449868
rect 3660 449828 3666 449840
rect 37918 449828 37924 449840
rect 37976 449828 37982 449880
rect 429102 448468 429108 448520
rect 429160 448508 429166 448520
rect 580902 448508 580908 448520
rect 429160 448480 580908 448508
rect 429160 448468 429166 448480
rect 580902 448468 580908 448480
rect 580960 448468 580966 448520
rect 6178 441532 6184 441584
rect 6236 441572 6242 441584
rect 37826 441572 37832 441584
rect 6236 441544 37832 441572
rect 6236 441532 6242 441544
rect 37826 441532 37832 441544
rect 37884 441532 37890 441584
rect 428642 438812 428648 438864
rect 428700 438852 428706 438864
rect 490558 438852 490564 438864
rect 428700 438824 490564 438852
rect 428700 438812 428706 438824
rect 490558 438812 490564 438824
rect 490616 438812 490622 438864
rect 3326 436092 3332 436144
rect 3384 436132 3390 436144
rect 11698 436132 11704 436144
rect 3384 436104 11704 436132
rect 3384 436092 3390 436104
rect 11698 436092 11704 436104
rect 11756 436092 11762 436144
rect 22738 431876 22744 431928
rect 22796 431916 22802 431928
rect 37826 431916 37832 431928
rect 22796 431888 37832 431916
rect 22796 431876 22802 431888
rect 37826 431876 37832 431888
rect 37884 431876 37890 431928
rect 428734 430584 428740 430636
rect 428792 430624 428798 430636
rect 580074 430624 580080 430636
rect 428792 430596 580080 430624
rect 428792 430584 428798 430596
rect 580074 430584 580080 430596
rect 580132 430584 580138 430636
rect 428642 429088 428648 429140
rect 428700 429128 428706 429140
rect 580258 429128 580264 429140
rect 428700 429100 580264 429128
rect 428700 429088 428706 429100
rect 580258 429088 580264 429100
rect 580316 429088 580322 429140
rect 3326 422288 3332 422340
rect 3384 422328 3390 422340
rect 26878 422328 26884 422340
rect 3384 422300 26884 422328
rect 3384 422288 3390 422300
rect 26878 422288 26884 422300
rect 26936 422288 26942 422340
rect 28258 422220 28264 422272
rect 28316 422260 28322 422272
rect 37918 422260 37924 422272
rect 28316 422232 37924 422260
rect 28316 422220 28322 422232
rect 37918 422220 37924 422232
rect 37976 422220 37982 422272
rect 428734 418140 428740 418192
rect 428792 418180 428798 418192
rect 580166 418180 580172 418192
rect 428792 418152 580172 418180
rect 428792 418140 428798 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3418 412564 3424 412616
rect 3476 412604 3482 412616
rect 37642 412604 37648 412616
rect 3476 412576 37648 412604
rect 3476 412564 3482 412576
rect 37642 412564 37648 412576
rect 37700 412564 37706 412616
rect 428826 409776 428832 409828
rect 428884 409816 428890 409828
rect 580350 409816 580356 409828
rect 428884 409788 580356 409816
rect 428884 409776 428890 409788
rect 580350 409776 580356 409788
rect 580408 409776 580414 409828
rect 3694 402908 3700 402960
rect 3752 402948 3758 402960
rect 37550 402948 37556 402960
rect 3752 402920 37556 402948
rect 3752 402908 3758 402920
rect 37550 402908 37556 402920
rect 37608 402908 37614 402960
rect 428458 400120 428464 400172
rect 428516 400160 428522 400172
rect 580442 400160 580448 400172
rect 428516 400132 580448 400160
rect 428516 400120 428522 400132
rect 580442 400120 580448 400132
rect 580500 400120 580506 400172
rect 10318 393252 10324 393304
rect 10376 393292 10382 393304
rect 37734 393292 37740 393304
rect 10376 393264 37740 393292
rect 10376 393252 10382 393264
rect 37734 393252 37740 393264
rect 37792 393252 37798 393304
rect 428458 390464 428464 390516
rect 428516 390504 428522 390516
rect 580534 390504 580540 390516
rect 428516 390476 580540 390504
rect 428516 390464 428522 390476
rect 580534 390464 580540 390476
rect 580592 390464 580598 390516
rect 3326 383664 3332 383716
rect 3384 383704 3390 383716
rect 24118 383704 24124 383716
rect 3384 383676 24124 383704
rect 3384 383664 3390 383676
rect 24118 383664 24124 383676
rect 24176 383664 24182 383716
rect 31018 383596 31024 383648
rect 31076 383636 31082 383648
rect 37458 383636 37464 383648
rect 31076 383608 37464 383636
rect 31076 383596 31082 383608
rect 37458 383596 37464 383608
rect 37516 383596 37522 383648
rect 3510 373940 3516 373992
rect 3568 373980 3574 373992
rect 37918 373980 37924 373992
rect 3568 373952 37924 373980
rect 3568 373940 3574 373952
rect 37918 373940 37924 373952
rect 37976 373940 37982 373992
rect 3142 371288 3148 371340
rect 3200 371328 3206 371340
rect 6178 371328 6184 371340
rect 3200 371300 6184 371328
rect 3200 371288 3206 371300
rect 6178 371288 6184 371300
rect 6236 371288 6242 371340
rect 428826 371152 428832 371204
rect 428884 371192 428890 371204
rect 580626 371192 580632 371204
rect 428884 371164 580632 371192
rect 428884 371152 428890 371164
rect 580626 371152 580632 371164
rect 580684 371152 580690 371204
rect 428458 364352 428464 364404
rect 428516 364392 428522 364404
rect 579798 364392 579804 364404
rect 428516 364364 579804 364392
rect 428516 364352 428522 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 3786 364284 3792 364336
rect 3844 364324 3850 364336
rect 37458 364324 37464 364336
rect 3844 364296 37464 364324
rect 3844 364284 3850 364296
rect 37458 364284 37464 364296
rect 37516 364284 37522 364336
rect 428550 361496 428556 361548
rect 428608 361536 428614 361548
rect 580718 361536 580724 361548
rect 428608 361508 580724 361536
rect 428608 361496 428614 361508
rect 580718 361496 580724 361508
rect 580776 361496 580782 361548
rect 11698 354628 11704 354680
rect 11756 354668 11762 354680
rect 37550 354668 37556 354680
rect 11756 354640 37556 354668
rect 11756 354628 11762 354640
rect 37550 354628 37556 354640
rect 37608 354628 37614 354680
rect 26878 344972 26884 345024
rect 26936 345012 26942 345024
rect 37642 345012 37648 345024
rect 26936 344984 37648 345012
rect 26936 344972 26942 344984
rect 37642 344972 37648 344984
rect 37700 344972 37706 345024
rect 3418 336676 3424 336728
rect 3476 336716 3482 336728
rect 37826 336716 37832 336728
rect 3476 336688 37832 336716
rect 3476 336676 3482 336688
rect 37826 336676 37832 336688
rect 37884 336676 37890 336728
rect 428550 332528 428556 332580
rect 428608 332568 428614 332580
rect 580258 332568 580264 332580
rect 428608 332540 580264 332568
rect 428608 332528 428614 332540
rect 580258 332528 580264 332540
rect 580316 332528 580322 332580
rect 2774 331576 2780 331628
rect 2832 331616 2838 331628
rect 4798 331616 4804 331628
rect 2832 331588 4804 331616
rect 2832 331576 2838 331588
rect 4798 331576 4804 331588
rect 4856 331576 4862 331628
rect 3602 327020 3608 327072
rect 3660 327060 3666 327072
rect 37550 327060 37556 327072
rect 3660 327032 37556 327060
rect 3660 327020 3666 327032
rect 37550 327020 37556 327032
rect 37608 327020 37614 327072
rect 428550 324300 428556 324352
rect 428608 324340 428614 324352
rect 579614 324340 579620 324352
rect 428608 324312 579620 324340
rect 428608 324300 428614 324312
rect 579614 324300 579620 324312
rect 579672 324300 579678 324352
rect 428826 322872 428832 322924
rect 428884 322912 428890 322924
rect 580350 322912 580356 322924
rect 428884 322884 580356 322912
rect 428884 322872 428890 322884
rect 580350 322872 580356 322884
rect 580408 322872 580414 322924
rect 24118 317364 24124 317416
rect 24176 317404 24182 317416
rect 37918 317404 37924 317416
rect 24176 317376 37924 317404
rect 24176 317364 24182 317376
rect 37918 317364 37924 317376
rect 37976 317364 37982 317416
rect 428734 313216 428740 313268
rect 428792 313256 428798 313268
rect 580442 313256 580448 313268
rect 428792 313228 580448 313256
rect 428792 313216 428798 313228
rect 580442 313216 580448 313228
rect 580500 313216 580506 313268
rect 428642 311856 428648 311908
rect 428700 311896 428706 311908
rect 580166 311896 580172 311908
rect 428700 311868 580172 311896
rect 428700 311856 428706 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 6178 307708 6184 307760
rect 6236 307748 6242 307760
rect 37366 307748 37372 307760
rect 6236 307720 37372 307748
rect 6236 307708 6242 307720
rect 37366 307708 37372 307720
rect 37424 307708 37430 307760
rect 3510 298052 3516 298104
rect 3568 298092 3574 298104
rect 37550 298092 37556 298104
rect 3568 298064 37556 298092
rect 3568 298052 3574 298064
rect 37550 298052 37556 298064
rect 37608 298052 37614 298104
rect 428458 292476 428464 292528
rect 428516 292516 428522 292528
rect 580534 292516 580540 292528
rect 428516 292488 580540 292516
rect 428516 292476 428522 292488
rect 580534 292476 580540 292488
rect 580592 292476 580598 292528
rect 3694 288328 3700 288380
rect 3752 288368 3758 288380
rect 37734 288368 37740 288380
rect 3752 288340 37740 288368
rect 3752 288328 3758 288340
rect 37734 288328 37740 288340
rect 37792 288328 37798 288380
rect 429010 282820 429016 282872
rect 429068 282860 429074 282872
rect 580626 282860 580632 282872
rect 429068 282832 580632 282860
rect 429068 282820 429074 282832
rect 580626 282820 580632 282832
rect 580684 282820 580690 282872
rect 4798 278672 4804 278724
rect 4856 278712 4862 278724
rect 37734 278712 37740 278724
rect 4856 278684 37740 278712
rect 4856 278672 4862 278684
rect 37734 278672 37740 278684
rect 37792 278672 37798 278724
rect 428458 271872 428464 271924
rect 428516 271912 428522 271924
rect 579614 271912 579620 271924
rect 428516 271884 579620 271912
rect 428516 271872 428522 271884
rect 579614 271872 579620 271884
rect 579672 271872 579678 271924
rect 3418 269016 3424 269068
rect 3476 269056 3482 269068
rect 37918 269056 37924 269068
rect 3476 269028 37924 269056
rect 3476 269016 3482 269028
rect 37918 269016 37924 269028
rect 37976 269016 37982 269068
rect 3602 259360 3608 259412
rect 3660 259400 3666 259412
rect 37366 259400 37372 259412
rect 3660 259372 37372 259400
rect 3660 259360 3666 259372
rect 37366 259360 37372 259372
rect 37424 259360 37430 259412
rect 428550 258068 428556 258120
rect 428608 258108 428614 258120
rect 579614 258108 579620 258120
rect 428608 258080 579620 258108
rect 428608 258068 428614 258080
rect 579614 258068 579620 258080
rect 579672 258068 579678 258120
rect 428918 253852 428924 253904
rect 428976 253892 428982 253904
rect 580258 253892 580264 253904
rect 428976 253864 580264 253892
rect 428976 253852 428982 253864
rect 580258 253852 580264 253864
rect 580316 253852 580322 253904
rect 3510 249704 3516 249756
rect 3568 249744 3574 249756
rect 37918 249744 37924 249756
rect 3568 249716 37924 249744
rect 3568 249704 3574 249716
rect 37918 249704 37924 249716
rect 37976 249704 37982 249756
rect 428734 244264 428740 244316
rect 428792 244304 428798 244316
rect 579798 244304 579804 244316
rect 428792 244276 579804 244304
rect 428792 244264 428798 244276
rect 579798 244264 579804 244276
rect 579856 244264 579862 244316
rect 428642 244196 428648 244248
rect 428700 244236 428706 244248
rect 580350 244236 580356 244248
rect 428700 244208 580356 244236
rect 428700 244196 428706 244208
rect 580350 244196 580356 244208
rect 580408 244196 580414 244248
rect 3694 240048 3700 240100
rect 3752 240088 3758 240100
rect 37366 240088 37372 240100
rect 3752 240060 37372 240088
rect 3752 240048 3758 240060
rect 37366 240048 37372 240060
rect 37424 240048 37430 240100
rect 428458 231820 428464 231872
rect 428516 231860 428522 231872
rect 580166 231860 580172 231872
rect 428516 231832 580172 231860
rect 428516 231820 428522 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 3418 231752 3424 231804
rect 3476 231792 3482 231804
rect 37642 231792 37648 231804
rect 3476 231764 37648 231792
rect 3476 231752 3482 231764
rect 37642 231752 37648 231764
rect 37700 231752 37706 231804
rect 3602 222096 3608 222148
rect 3660 222136 3666 222148
rect 37734 222136 37740 222148
rect 3660 222108 37740 222136
rect 3660 222096 3666 222108
rect 37734 222096 37740 222108
rect 37792 222096 37798 222148
rect 428550 218016 428556 218068
rect 428608 218056 428614 218068
rect 580166 218056 580172 218068
rect 428608 218028 580172 218056
rect 428608 218016 428614 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 3510 212440 3516 212492
rect 3568 212480 3574 212492
rect 37826 212480 37832 212492
rect 3568 212452 37832 212480
rect 3568 212440 3574 212452
rect 37826 212440 37832 212452
rect 37884 212440 37890 212492
rect 428642 205640 428648 205692
rect 428700 205680 428706 205692
rect 580166 205680 580172 205692
rect 428700 205652 580172 205680
rect 428700 205640 428706 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 37734 202824 37740 202836
rect 3476 202796 37740 202824
rect 3476 202784 3482 202796
rect 37734 202784 37740 202796
rect 37792 202784 37798 202836
rect 3602 193128 3608 193180
rect 3660 193168 3666 193180
rect 37734 193168 37740 193180
rect 3660 193140 37740 193168
rect 3660 193128 3666 193140
rect 37734 193128 37740 193140
rect 37792 193128 37798 193180
rect 428458 191836 428464 191888
rect 428516 191876 428522 191888
rect 580166 191876 580172 191888
rect 428516 191848 580172 191876
rect 428516 191836 428522 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 3510 183472 3516 183524
rect 3568 183512 3574 183524
rect 37918 183512 37924 183524
rect 3568 183484 37924 183512
rect 3568 183472 3574 183484
rect 37918 183472 37924 183484
rect 37976 183472 37982 183524
rect 428550 178032 428556 178084
rect 428608 178072 428614 178084
rect 580166 178072 580172 178084
rect 428608 178044 580172 178072
rect 428608 178032 428614 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 3418 173816 3424 173868
rect 3476 173856 3482 173868
rect 37734 173856 37740 173868
rect 3476 173828 37740 173856
rect 3476 173816 3482 173828
rect 37734 173816 37740 173828
rect 37792 173816 37798 173868
rect 428458 165588 428464 165640
rect 428516 165628 428522 165640
rect 580166 165628 580172 165640
rect 428516 165600 580172 165628
rect 428516 165588 428522 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 3510 164160 3516 164212
rect 3568 164200 3574 164212
rect 37918 164200 37924 164212
rect 3568 164172 37924 164200
rect 3568 164160 3574 164172
rect 37918 164160 37924 164172
rect 37976 164160 37982 164212
rect 3418 154504 3424 154556
rect 3476 154544 3482 154556
rect 37642 154544 37648 154556
rect 3476 154516 37648 154544
rect 3476 154504 3482 154516
rect 37642 154504 37648 154516
rect 37700 154504 37706 154556
rect 429102 151784 429108 151836
rect 429160 151824 429166 151836
rect 579982 151824 579988 151836
rect 429160 151796 579988 151824
rect 429160 151784 429166 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3326 144848 3332 144900
rect 3384 144888 3390 144900
rect 37918 144888 37924 144900
rect 3384 144860 37924 144888
rect 3384 144848 3390 144860
rect 37918 144848 37924 144860
rect 37976 144848 37982 144900
rect 428826 137980 428832 138032
rect 428884 138020 428890 138032
rect 580166 138020 580172 138032
rect 428884 137992 580172 138020
rect 428884 137980 428890 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 3418 136552 3424 136604
rect 3476 136592 3482 136604
rect 37550 136592 37556 136604
rect 3476 136564 37556 136592
rect 3476 136552 3482 136564
rect 37550 136552 37556 136564
rect 37608 136552 37614 136604
rect 428918 126896 428924 126948
rect 428976 126936 428982 126948
rect 580166 126936 580172 126948
rect 428976 126908 580172 126936
rect 428976 126896 428982 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3418 124108 3424 124160
rect 3476 124148 3482 124160
rect 37734 124148 37740 124160
rect 3476 124120 37740 124148
rect 3476 124108 3482 124120
rect 37734 124108 37740 124120
rect 37792 124108 37798 124160
rect 428458 113092 428464 113144
rect 428516 113132 428522 113144
rect 579798 113132 579804 113144
rect 428516 113104 579804 113132
rect 428516 113092 428522 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 37918 111772 37924 111784
rect 3476 111744 37924 111772
rect 3476 111732 3482 111744
rect 37918 111732 37924 111744
rect 37976 111732 37982 111784
rect 428458 100648 428464 100700
rect 428516 100688 428522 100700
rect 580166 100688 580172 100700
rect 428516 100660 580172 100688
rect 428516 100648 428522 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 37918 97968 37924 97980
rect 3476 97940 37924 97968
rect 3476 97928 3482 97940
rect 37918 97928 37924 97940
rect 37976 97928 37982 97980
rect 428550 86912 428556 86964
rect 428608 86952 428614 86964
rect 580166 86952 580172 86964
rect 428608 86924 580172 86952
rect 428608 86912 428614 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 38010 85524 38016 85536
rect 3200 85496 38016 85524
rect 3200 85484 3206 85496
rect 38010 85484 38016 85496
rect 38068 85484 38074 85536
rect 428458 73108 428464 73160
rect 428516 73148 428522 73160
rect 580166 73148 580172 73160
rect 428516 73120 580172 73148
rect 428516 73108 428522 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 37918 71720 37924 71732
rect 3476 71692 37924 71720
rect 3476 71680 3482 71692
rect 37918 71680 37924 71692
rect 37976 71680 37982 71732
rect 428550 60664 428556 60716
rect 428608 60704 428614 60716
rect 580166 60704 580172 60716
rect 428608 60676 580172 60704
rect 428608 60664 428614 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 38010 59344 38016 59356
rect 3108 59316 38016 59344
rect 3108 59304 3114 59316
rect 38010 59304 38016 59316
rect 38068 59304 38074 59356
rect 428458 46860 428464 46912
rect 428516 46900 428522 46912
rect 580166 46900 580172 46912
rect 428516 46872 580172 46900
rect 428516 46860 428522 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 37918 45540 37924 45552
rect 3476 45512 37924 45540
rect 3476 45500 3482 45512
rect 37918 45500 37924 45512
rect 37976 45500 37982 45552
rect 212534 39516 212540 39568
rect 212592 39556 212598 39568
rect 212902 39556 212908 39568
rect 212592 39528 212908 39556
rect 212592 39516 212598 39528
rect 212902 39516 212908 39528
rect 212960 39516 212966 39568
rect 72418 38564 72424 38616
rect 72476 38604 72482 38616
rect 73982 38604 73988 38616
rect 72476 38576 73988 38604
rect 72476 38564 72482 38576
rect 73982 38564 73988 38576
rect 74040 38564 74046 38616
rect 194042 38428 194048 38480
rect 194100 38468 194106 38480
rect 195238 38468 195244 38480
rect 194100 38440 195244 38468
rect 194100 38428 194106 38440
rect 195238 38428 195244 38440
rect 195296 38428 195302 38480
rect 297082 38428 297088 38480
rect 297140 38468 297146 38480
rect 312538 38468 312544 38480
rect 297140 38440 312544 38468
rect 297140 38428 297146 38440
rect 312538 38428 312544 38440
rect 312596 38428 312602 38480
rect 55858 38360 55864 38412
rect 55916 38400 55922 38412
rect 58618 38400 58624 38412
rect 55916 38372 58624 38400
rect 55916 38360 55922 38372
rect 58618 38360 58624 38372
rect 58676 38360 58682 38412
rect 207290 38360 207296 38412
rect 207348 38400 207354 38412
rect 209038 38400 209044 38412
rect 207348 38372 209044 38400
rect 207348 38360 207354 38372
rect 209038 38360 209044 38372
rect 209096 38360 209102 38412
rect 311802 38360 311808 38412
rect 311860 38400 311866 38412
rect 349798 38400 349804 38412
rect 311860 38372 349804 38400
rect 311860 38360 311866 38372
rect 349798 38360 349804 38372
rect 349856 38360 349862 38412
rect 47578 38292 47584 38344
rect 47636 38332 47642 38344
rect 48314 38332 48320 38344
rect 47636 38304 48320 38332
rect 47636 38292 47642 38304
rect 48314 38292 48320 38304
rect 48372 38292 48378 38344
rect 282178 38292 282184 38344
rect 282236 38332 282242 38344
rect 324590 38332 324596 38344
rect 282236 38304 324596 38332
rect 282236 38292 282242 38304
rect 324590 38292 324596 38304
rect 324648 38292 324654 38344
rect 324958 38292 324964 38344
rect 325016 38332 325022 38344
rect 356606 38332 356612 38344
rect 325016 38304 356612 38332
rect 325016 38292 325022 38304
rect 356606 38292 356612 38304
rect 356664 38292 356670 38344
rect 411806 38292 411812 38344
rect 411864 38332 411870 38344
rect 425698 38332 425704 38344
rect 411864 38304 425704 38332
rect 411864 38292 411870 38304
rect 425698 38292 425704 38304
rect 425756 38292 425762 38344
rect 46198 38224 46204 38276
rect 46256 38264 46262 38276
rect 48958 38264 48964 38276
rect 46256 38236 48964 38264
rect 46256 38224 46262 38236
rect 48958 38224 48964 38236
rect 49016 38224 49022 38276
rect 185394 38224 185400 38276
rect 185452 38264 185458 38276
rect 188338 38264 188344 38276
rect 185452 38236 188344 38264
rect 185452 38224 185458 38236
rect 188338 38224 188344 38236
rect 188396 38224 188402 38276
rect 203426 38224 203432 38276
rect 203484 38264 203490 38276
rect 224126 38264 224132 38276
rect 203484 38236 224132 38264
rect 203484 38224 203490 38236
rect 224126 38224 224132 38236
rect 224184 38224 224190 38276
rect 286318 38224 286324 38276
rect 286376 38264 286382 38276
rect 330018 38264 330024 38276
rect 286376 38236 330024 38264
rect 286376 38224 286382 38236
rect 330018 38224 330024 38236
rect 330076 38224 330082 38276
rect 330570 38224 330576 38276
rect 330628 38264 330634 38276
rect 348786 38264 348792 38276
rect 330628 38236 348792 38264
rect 330628 38224 330634 38236
rect 348786 38224 348792 38236
rect 348844 38224 348850 38276
rect 375374 38224 375380 38276
rect 375432 38264 375438 38276
rect 376846 38264 376852 38276
rect 375432 38236 376852 38264
rect 375432 38224 375438 38236
rect 376846 38224 376852 38236
rect 376904 38224 376910 38276
rect 393038 38224 393044 38276
rect 393096 38264 393102 38276
rect 447134 38264 447140 38276
rect 393096 38236 447140 38264
rect 393096 38224 393102 38236
rect 447134 38224 447140 38236
rect 447192 38224 447198 38276
rect 75914 38156 75920 38208
rect 75972 38196 75978 38208
rect 77294 38196 77300 38208
rect 75972 38168 77300 38196
rect 75972 38156 75978 38168
rect 77294 38156 77300 38168
rect 77352 38156 77358 38208
rect 163590 38156 163596 38208
rect 163648 38196 163654 38208
rect 170398 38196 170404 38208
rect 163648 38168 170404 38196
rect 163648 38156 163654 38168
rect 170398 38156 170404 38168
rect 170456 38156 170462 38208
rect 171318 38156 171324 38208
rect 171376 38196 171382 38208
rect 172698 38196 172704 38208
rect 171376 38168 172704 38196
rect 171376 38156 171382 38168
rect 172698 38156 172704 38168
rect 172756 38156 172762 38208
rect 181530 38156 181536 38208
rect 181588 38196 181594 38208
rect 218698 38196 218704 38208
rect 181588 38168 218704 38196
rect 181588 38156 181594 38168
rect 218698 38156 218704 38168
rect 218756 38156 218762 38208
rect 226610 38156 226616 38208
rect 226668 38196 226674 38208
rect 244274 38196 244280 38208
rect 226668 38168 244280 38196
rect 226668 38156 226674 38168
rect 244274 38156 244280 38168
rect 244332 38156 244338 38208
rect 277210 38156 277216 38208
rect 277268 38196 277274 38208
rect 307110 38196 307116 38208
rect 277268 38168 307116 38196
rect 277268 38156 277274 38168
rect 307110 38156 307116 38168
rect 307168 38156 307174 38208
rect 322014 38156 322020 38208
rect 322072 38196 322078 38208
rect 414658 38196 414664 38208
rect 322072 38168 414664 38196
rect 322072 38156 322078 38168
rect 414658 38156 414664 38168
rect 414716 38156 414722 38208
rect 415670 38156 415676 38208
rect 415728 38196 415734 38208
rect 436738 38196 436744 38208
rect 415728 38168 436744 38196
rect 415728 38156 415734 38168
rect 436738 38156 436744 38168
rect 436796 38156 436802 38208
rect 66806 38088 66812 38140
rect 66864 38128 66870 38140
rect 68922 38128 68928 38140
rect 66864 38100 68928 38128
rect 66864 38088 66870 38100
rect 68922 38088 68928 38100
rect 68980 38088 68986 38140
rect 169662 38088 169668 38140
rect 169720 38128 169726 38140
rect 200758 38128 200764 38140
rect 169720 38100 200764 38128
rect 169720 38088 169726 38100
rect 200758 38088 200764 38100
rect 200816 38088 200822 38140
rect 215846 38088 215852 38140
rect 215904 38128 215910 38140
rect 342898 38128 342904 38140
rect 215904 38100 342904 38128
rect 215904 38088 215910 38100
rect 342898 38088 342904 38100
rect 342956 38088 342962 38140
rect 394602 38088 394608 38140
rect 394660 38128 394666 38140
rect 454034 38128 454040 38140
rect 394660 38100 454040 38128
rect 394660 38088 394666 38100
rect 454034 38088 454040 38100
rect 454092 38088 454098 38140
rect 59722 38020 59728 38072
rect 59780 38060 59786 38072
rect 69658 38060 69664 38072
rect 59780 38032 69664 38060
rect 59780 38020 59786 38032
rect 69658 38020 69664 38032
rect 69716 38020 69722 38072
rect 84746 38020 84752 38072
rect 84804 38060 84810 38072
rect 86954 38060 86960 38072
rect 84804 38032 86960 38060
rect 84804 38020 84810 38032
rect 86954 38020 86960 38032
rect 87012 38020 87018 38072
rect 91002 38020 91008 38072
rect 91060 38060 91066 38072
rect 93118 38060 93124 38072
rect 91060 38032 93124 38060
rect 91060 38020 91066 38032
rect 93118 38020 93124 38032
rect 93176 38020 93182 38072
rect 97994 38020 98000 38072
rect 98052 38060 98058 38072
rect 99006 38060 99012 38072
rect 98052 38032 99012 38060
rect 98052 38020 98058 38032
rect 99006 38020 99012 38032
rect 99064 38020 99070 38072
rect 101398 38020 101404 38072
rect 101456 38060 101462 38072
rect 102134 38060 102140 38072
rect 101456 38032 102140 38060
rect 101456 38020 101462 38032
rect 102134 38020 102140 38032
rect 102192 38020 102198 38072
rect 105538 38060 105544 38072
rect 103486 38032 105544 38060
rect 39298 37952 39304 38004
rect 39356 37992 39362 38004
rect 40494 37992 40500 38004
rect 39356 37964 40500 37992
rect 39356 37952 39362 37964
rect 40494 37952 40500 37964
rect 40552 37952 40558 38004
rect 41322 37952 41328 38004
rect 41380 37992 41386 38004
rect 41966 37992 41972 38004
rect 41380 37964 41972 37992
rect 41380 37952 41386 37964
rect 41966 37952 41972 37964
rect 42024 37952 42030 38004
rect 44174 37952 44180 38004
rect 44232 37992 44238 38004
rect 45094 37992 45100 38004
rect 44232 37964 45100 37992
rect 44232 37952 44238 37964
rect 45094 37952 45100 37964
rect 45152 37952 45158 38004
rect 49694 37952 49700 38004
rect 49752 37992 49758 38004
rect 50614 37992 50620 38004
rect 49752 37964 50620 37992
rect 49752 37952 49758 37964
rect 50614 37952 50620 37964
rect 50672 37952 50678 38004
rect 52454 37952 52460 38004
rect 52512 37992 52518 38004
rect 52914 37992 52920 38004
rect 52512 37964 52920 37992
rect 52512 37952 52518 37964
rect 52914 37952 52920 37964
rect 52972 37952 52978 38004
rect 56594 37952 56600 38004
rect 56652 37992 56658 38004
rect 57606 37992 57612 38004
rect 56652 37964 57612 37992
rect 56652 37952 56658 37964
rect 57606 37952 57612 37964
rect 57664 37952 57670 38004
rect 62114 37952 62120 38004
rect 62172 37992 62178 38004
rect 63126 37992 63132 38004
rect 62172 37964 63132 37992
rect 62172 37952 62178 37964
rect 63126 37952 63132 37964
rect 63184 37952 63190 38004
rect 64874 37952 64880 38004
rect 64932 37992 64938 38004
rect 65426 37992 65432 38004
rect 64932 37964 65432 37992
rect 64932 37952 64938 37964
rect 65426 37952 65432 37964
rect 65484 37952 65490 38004
rect 70394 37952 70400 38004
rect 70452 37992 70458 38004
rect 70854 37992 70860 38004
rect 70452 37964 70860 37992
rect 70452 37952 70458 37964
rect 70854 37952 70860 37964
rect 70912 37952 70918 38004
rect 71038 37952 71044 38004
rect 71096 37992 71102 38004
rect 73246 37992 73252 38004
rect 71096 37964 73252 37992
rect 71096 37952 71102 37964
rect 73246 37952 73252 37964
rect 73304 37952 73310 38004
rect 74534 37952 74540 38004
rect 74592 37992 74598 38004
rect 75546 37992 75552 38004
rect 74592 37964 75552 37992
rect 74592 37952 74598 37964
rect 75546 37952 75552 37964
rect 75604 37952 75610 38004
rect 80054 37952 80060 38004
rect 80112 37992 80118 38004
rect 80974 37992 80980 38004
rect 80112 37964 80980 37992
rect 80112 37952 80118 37964
rect 80974 37952 80980 37964
rect 81032 37952 81038 38004
rect 85574 37952 85580 38004
rect 85632 37992 85638 38004
rect 86494 37992 86500 38004
rect 85632 37964 86500 37992
rect 85632 37952 85638 37964
rect 86494 37952 86500 37964
rect 86552 37952 86558 38004
rect 88334 37952 88340 38004
rect 88392 37992 88398 38004
rect 88886 37992 88892 38004
rect 88392 37964 88892 37992
rect 88392 37952 88398 37964
rect 88886 37952 88892 37964
rect 88944 37952 88950 38004
rect 91738 37952 91744 38004
rect 91796 37992 91802 38004
rect 103486 37992 103514 38032
rect 105538 38020 105544 38032
rect 105596 38020 105602 38072
rect 130746 38020 130752 38072
rect 130804 38060 130810 38072
rect 141418 38060 141424 38072
rect 130804 38032 141424 38060
rect 130804 38020 130810 38032
rect 141418 38020 141424 38032
rect 141476 38020 141482 38072
rect 142154 38020 142160 38072
rect 142212 38060 142218 38072
rect 142614 38060 142620 38072
rect 142212 38032 142620 38060
rect 142212 38020 142218 38032
rect 142614 38020 142620 38032
rect 142672 38020 142678 38072
rect 154666 38020 154672 38072
rect 154724 38060 154730 38072
rect 155126 38060 155132 38072
rect 154724 38032 155132 38060
rect 154724 38020 154730 38032
rect 155126 38020 155132 38032
rect 155184 38020 155190 38072
rect 165614 38020 165620 38072
rect 165672 38060 165678 38072
rect 166166 38060 166172 38072
rect 165672 38032 166172 38060
rect 165672 38020 165678 38032
rect 166166 38020 166172 38032
rect 166224 38020 166230 38072
rect 199470 38020 199476 38072
rect 199528 38060 199534 38072
rect 328730 38060 328736 38072
rect 199528 38032 328736 38060
rect 199528 38020 199534 38032
rect 328730 38020 328736 38032
rect 328788 38020 328794 38072
rect 330478 38020 330484 38072
rect 330536 38060 330542 38072
rect 332594 38060 332600 38072
rect 330536 38032 332600 38060
rect 330536 38020 330542 38032
rect 332594 38020 332600 38032
rect 332652 38020 332658 38072
rect 335354 38020 335360 38072
rect 335412 38060 335418 38072
rect 336274 38060 336280 38072
rect 335412 38032 336280 38060
rect 335412 38020 335418 38032
rect 336274 38020 336280 38032
rect 336332 38020 336338 38072
rect 340138 38020 340144 38072
rect 340196 38060 340202 38072
rect 340874 38060 340880 38072
rect 340196 38032 340880 38060
rect 340196 38020 340202 38032
rect 340874 38020 340880 38032
rect 340932 38020 340938 38072
rect 341058 38020 341064 38072
rect 341116 38060 341122 38072
rect 369118 38060 369124 38072
rect 341116 38032 369124 38060
rect 341116 38020 341122 38032
rect 369118 38020 369124 38032
rect 369176 38020 369182 38072
rect 382826 38020 382832 38072
rect 382884 38060 382890 38072
rect 392578 38060 392584 38072
rect 382884 38032 392584 38060
rect 382884 38020 382890 38032
rect 392578 38020 392584 38032
rect 392636 38020 392642 38072
rect 395890 38020 395896 38072
rect 395948 38060 395954 38072
rect 460934 38060 460940 38072
rect 395948 38032 460940 38060
rect 395948 38020 395954 38032
rect 460934 38020 460940 38032
rect 460992 38020 460998 38072
rect 91796 37964 103514 37992
rect 91796 37952 91802 37964
rect 104158 37952 104164 38004
rect 104216 37992 104222 38004
rect 106274 37992 106280 38004
rect 104216 37964 106280 37992
rect 104216 37952 104222 37964
rect 106274 37952 106280 37964
rect 106332 37952 106338 38004
rect 115842 37952 115848 38004
rect 115900 37992 115906 38004
rect 116578 37992 116584 38004
rect 115900 37964 116584 37992
rect 115900 37952 115906 37964
rect 116578 37952 116584 37964
rect 116636 37952 116642 38004
rect 124214 37952 124220 38004
rect 124272 37992 124278 38004
rect 124766 37992 124772 38004
rect 124272 37964 124772 37992
rect 124272 37952 124278 37964
rect 124766 37952 124772 37964
rect 124824 37952 124830 38004
rect 128262 37952 128268 38004
rect 128320 37992 128326 38004
rect 128998 37992 129004 38004
rect 128320 37964 129004 37992
rect 128320 37952 128326 37964
rect 128998 37952 129004 37964
rect 129056 37952 129062 38004
rect 132126 37952 132132 38004
rect 132184 37992 132190 38004
rect 146938 37992 146944 38004
rect 132184 37964 146944 37992
rect 132184 37952 132190 37964
rect 146938 37952 146944 37964
rect 146996 37952 147002 38004
rect 148778 37952 148784 38004
rect 148836 37992 148842 38004
rect 217318 37992 217324 38004
rect 148836 37964 217324 37992
rect 148836 37952 148842 37964
rect 217318 37952 217324 37964
rect 217376 37952 217382 38004
rect 218790 37952 218796 38004
rect 218848 37992 218854 38004
rect 218848 37964 356560 37992
rect 218848 37952 218854 37964
rect 10318 37884 10324 37936
rect 10376 37924 10382 37936
rect 121638 37924 121644 37936
rect 10376 37896 121644 37924
rect 10376 37884 10382 37896
rect 121638 37884 121644 37896
rect 121696 37884 121702 37936
rect 136266 37884 136272 37936
rect 136324 37924 136330 37936
rect 177298 37924 177304 37936
rect 136324 37896 177304 37924
rect 136324 37884 136330 37896
rect 177298 37884 177304 37896
rect 177356 37884 177362 37936
rect 186958 37884 186964 37936
rect 187016 37924 187022 37936
rect 187016 37896 354674 37924
rect 187016 37884 187022 37896
rect 75178 37816 75184 37868
rect 75236 37856 75242 37868
rect 77846 37856 77852 37868
rect 75236 37828 77852 37856
rect 75236 37816 75242 37828
rect 77846 37816 77852 37828
rect 77904 37816 77910 37868
rect 149514 37816 149520 37868
rect 149572 37856 149578 37868
rect 150618 37856 150624 37868
rect 149572 37828 150624 37856
rect 149572 37816 149578 37828
rect 150618 37816 150624 37828
rect 150676 37816 150682 37868
rect 204162 37816 204168 37868
rect 204220 37856 204226 37868
rect 206922 37856 206928 37868
rect 204220 37828 206928 37856
rect 204220 37816 204226 37828
rect 206922 37816 206928 37828
rect 206980 37816 206986 37868
rect 219434 37816 219440 37868
rect 219492 37856 219498 37868
rect 219986 37856 219992 37868
rect 219492 37828 219992 37856
rect 219492 37816 219498 37828
rect 219986 37816 219992 37828
rect 220044 37816 220050 37868
rect 222102 37816 222108 37868
rect 222160 37856 222166 37868
rect 222654 37856 222660 37868
rect 222160 37828 222660 37856
rect 222160 37816 222166 37828
rect 222654 37816 222660 37828
rect 222712 37816 222718 37868
rect 224218 37816 224224 37868
rect 224276 37856 224282 37868
rect 224954 37856 224960 37868
rect 224276 37828 224960 37856
rect 224276 37816 224282 37828
rect 224954 37816 224960 37828
rect 225012 37816 225018 37868
rect 242158 37816 242164 37868
rect 242216 37856 242222 37868
rect 242894 37856 242900 37868
rect 242216 37828 242900 37856
rect 242216 37816 242222 37828
rect 242894 37816 242900 37828
rect 242952 37816 242958 37868
rect 244918 37816 244924 37868
rect 244976 37856 244982 37868
rect 245746 37856 245752 37868
rect 244976 37828 245752 37856
rect 244976 37816 244982 37828
rect 245746 37816 245752 37828
rect 245804 37816 245810 37868
rect 248414 37816 248420 37868
rect 248472 37856 248478 37868
rect 248874 37856 248880 37868
rect 248472 37828 248880 37856
rect 248472 37816 248478 37828
rect 248874 37816 248880 37828
rect 248932 37816 248938 37868
rect 252554 37816 252560 37868
rect 252612 37856 252618 37868
rect 253566 37856 253572 37868
rect 252612 37828 253572 37856
rect 252612 37816 252618 37828
rect 253566 37816 253572 37828
rect 253624 37816 253630 37868
rect 261110 37816 261116 37868
rect 261168 37856 261174 37868
rect 262858 37856 262864 37868
rect 261168 37828 262864 37856
rect 261168 37816 261174 37828
rect 262858 37816 262864 37828
rect 262916 37816 262922 37868
rect 266354 37816 266360 37868
rect 266412 37856 266418 37868
rect 266814 37856 266820 37868
rect 266412 37828 266820 37856
rect 266412 37816 266418 37828
rect 266814 37816 266820 37828
rect 266872 37816 266878 37868
rect 284294 37816 284300 37868
rect 284352 37856 284358 37868
rect 284754 37856 284760 37868
rect 284352 37828 284760 37856
rect 284352 37816 284358 37828
rect 284754 37816 284760 37828
rect 284812 37816 284818 37868
rect 288434 37816 288440 37868
rect 288492 37856 288498 37868
rect 289446 37856 289452 37868
rect 288492 37828 289452 37856
rect 288492 37816 288498 37828
rect 289446 37816 289452 37828
rect 289504 37816 289510 37868
rect 294046 37816 294052 37868
rect 294104 37856 294110 37868
rect 294966 37856 294972 37868
rect 294104 37828 294972 37856
rect 294104 37816 294110 37828
rect 294966 37816 294972 37828
rect 295024 37816 295030 37868
rect 308030 37816 308036 37868
rect 308088 37856 308094 37868
rect 309778 37856 309784 37868
rect 308088 37828 309784 37856
rect 308088 37816 308094 37828
rect 309778 37816 309784 37828
rect 309836 37816 309842 37868
rect 320174 37816 320180 37868
rect 320232 37856 320238 37868
rect 320726 37856 320732 37868
rect 320232 37828 320732 37856
rect 320232 37816 320238 37828
rect 320726 37816 320732 37828
rect 320784 37816 320790 37868
rect 322198 37816 322204 37868
rect 322256 37856 322262 37868
rect 323026 37856 323032 37868
rect 322256 37828 323032 37856
rect 322256 37816 322262 37828
rect 323026 37816 323032 37828
rect 323084 37816 323090 37868
rect 325694 37816 325700 37868
rect 325752 37856 325758 37868
rect 326154 37856 326160 37868
rect 325752 37828 326160 37856
rect 325752 37816 325758 37828
rect 326154 37816 326160 37828
rect 326212 37816 326218 37868
rect 328730 37816 328736 37868
rect 328788 37856 328794 37868
rect 331858 37856 331864 37868
rect 328788 37828 331864 37856
rect 328788 37816 328794 37828
rect 331858 37816 331864 37828
rect 331916 37816 331922 37868
rect 348418 37816 348424 37868
rect 348476 37856 348482 37868
rect 350534 37856 350540 37868
rect 348476 37828 350540 37856
rect 348476 37816 348482 37828
rect 350534 37816 350540 37828
rect 350592 37816 350598 37868
rect 293126 37748 293132 37800
rect 293184 37788 293190 37800
rect 295978 37788 295984 37800
rect 293184 37760 295984 37788
rect 293184 37748 293190 37760
rect 295978 37748 295984 37760
rect 296036 37748 296042 37800
rect 354646 37788 354674 37896
rect 356532 37856 356560 37964
rect 356698 37952 356704 38004
rect 356756 37992 356762 38004
rect 358906 37992 358912 38004
rect 356756 37964 358912 37992
rect 356756 37952 356762 37964
rect 358906 37952 358912 37964
rect 358964 37952 358970 38004
rect 365714 37952 365720 38004
rect 365772 37992 365778 38004
rect 366726 37992 366732 38004
rect 365772 37964 366732 37992
rect 365772 37952 365778 37964
rect 366726 37952 366732 37964
rect 366784 37952 366790 38004
rect 385034 37952 385040 38004
rect 385092 37992 385098 38004
rect 385494 37992 385500 38004
rect 385092 37964 385500 37992
rect 385092 37952 385098 37964
rect 385494 37952 385500 37964
rect 385552 37952 385558 38004
rect 389174 37952 389180 38004
rect 389232 37992 389238 38004
rect 390094 37992 390100 38004
rect 389232 37964 390100 37992
rect 389232 37952 389238 37964
rect 390094 37952 390100 37964
rect 390152 37952 390158 38004
rect 397730 37952 397736 38004
rect 397788 37992 397794 38004
rect 467834 37992 467840 38004
rect 397788 37964 467840 37992
rect 397788 37952 397794 37964
rect 467834 37952 467840 37964
rect 467892 37952 467898 38004
rect 393958 37924 393964 37936
rect 364306 37896 393964 37924
rect 360838 37856 360844 37868
rect 356532 37828 360844 37856
rect 360838 37816 360844 37828
rect 360896 37816 360902 37868
rect 364306 37788 364334 37896
rect 393958 37884 393964 37896
rect 394016 37884 394022 37936
rect 399294 37884 399300 37936
rect 399352 37924 399358 37936
rect 474734 37924 474740 37936
rect 399352 37896 474740 37924
rect 399352 37884 399358 37896
rect 474734 37884 474740 37896
rect 474792 37884 474798 37936
rect 420914 37816 420920 37868
rect 420972 37856 420978 37868
rect 421374 37856 421380 37868
rect 420972 37828 421380 37856
rect 420972 37816 420978 37828
rect 421374 37816 421380 37828
rect 421432 37816 421438 37868
rect 354646 37760 364334 37788
rect 131574 37612 131580 37664
rect 131632 37652 131638 37664
rect 133782 37652 133788 37664
rect 131632 37624 133788 37652
rect 131632 37612 131638 37624
rect 133782 37612 133788 37624
rect 133840 37612 133846 37664
rect 189166 37612 189172 37664
rect 189224 37652 189230 37664
rect 190638 37652 190644 37664
rect 189224 37624 190644 37652
rect 189224 37612 189230 37624
rect 190638 37612 190644 37624
rect 190696 37612 190702 37664
rect 279050 37612 279056 37664
rect 279108 37652 279114 37664
rect 280798 37652 280804 37664
rect 279108 37624 280804 37652
rect 279108 37612 279114 37624
rect 280798 37612 280804 37624
rect 280856 37612 280862 37664
rect 106274 37340 106280 37392
rect 106332 37380 106338 37392
rect 113266 37380 113272 37392
rect 106332 37352 113272 37380
rect 106332 37340 106338 37352
rect 113266 37340 113272 37352
rect 113324 37340 113330 37392
rect 110414 37272 110420 37324
rect 110472 37312 110478 37324
rect 114002 37312 114008 37324
rect 110472 37284 114008 37312
rect 110472 37272 110478 37284
rect 114002 37272 114008 37284
rect 114060 37272 114066 37324
rect 275186 37272 275192 37324
rect 275244 37312 275250 37324
rect 275244 37284 277440 37312
rect 275244 37272 275250 37284
rect 277412 37244 277440 37284
rect 315022 37272 315028 37324
rect 315080 37312 315086 37324
rect 318058 37312 318064 37324
rect 315080 37284 318064 37312
rect 315080 37272 315086 37284
rect 318058 37272 318064 37284
rect 318116 37272 318122 37324
rect 353938 37272 353944 37324
rect 353996 37312 354002 37324
rect 355042 37312 355048 37324
rect 353996 37284 355048 37312
rect 353996 37272 354002 37284
rect 355042 37272 355048 37284
rect 355100 37272 355106 37324
rect 277412 37216 282914 37244
rect 282886 36972 282914 37216
rect 364334 36972 364340 36984
rect 282886 36944 364340 36972
rect 364334 36932 364340 36944
rect 364392 36932 364398 36984
rect 223574 36864 223580 36916
rect 223632 36904 223638 36916
rect 343542 36904 343548 36916
rect 223632 36876 343548 36904
rect 223632 36864 223638 36876
rect 343542 36864 343548 36876
rect 343600 36864 343606 36916
rect 167454 36796 167460 36848
rect 167512 36836 167518 36848
rect 327074 36836 327080 36848
rect 167512 36808 327080 36836
rect 167512 36796 167518 36808
rect 327074 36796 327080 36808
rect 327132 36796 327138 36848
rect 154574 36728 154580 36780
rect 154632 36768 154638 36780
rect 228542 36768 228548 36780
rect 154632 36740 228548 36768
rect 154632 36728 154638 36740
rect 228542 36728 228548 36740
rect 228600 36728 228606 36780
rect 297818 36728 297824 36780
rect 297876 36768 297882 36780
rect 466454 36768 466460 36780
rect 297876 36740 466460 36768
rect 297876 36728 297882 36740
rect 466454 36728 466460 36740
rect 466512 36728 466518 36780
rect 156506 36660 156512 36712
rect 156564 36700 156570 36712
rect 277394 36700 277400 36712
rect 156564 36672 277400 36700
rect 156564 36660 156570 36672
rect 277394 36660 277400 36672
rect 277452 36660 277458 36712
rect 313182 36660 313188 36712
rect 313240 36700 313246 36712
rect 538214 36700 538220 36712
rect 313240 36672 538220 36700
rect 313240 36660 313246 36672
rect 538214 36660 538220 36672
rect 538272 36660 538278 36712
rect 4798 36592 4804 36644
rect 4856 36632 4862 36644
rect 41414 36632 41420 36644
rect 4856 36604 41420 36632
rect 4856 36592 4862 36604
rect 41414 36592 41420 36604
rect 41472 36592 41478 36644
rect 56502 36592 56508 36644
rect 56560 36632 56566 36644
rect 76098 36632 76104 36644
rect 56560 36604 76104 36632
rect 56560 36592 56566 36604
rect 76098 36592 76104 36604
rect 76156 36592 76162 36644
rect 92382 36592 92388 36644
rect 92440 36632 92446 36644
rect 122834 36632 122840 36644
rect 92440 36604 122840 36632
rect 92440 36592 92446 36604
rect 122834 36592 122840 36604
rect 122892 36592 122898 36644
rect 217870 36592 217876 36644
rect 217928 36632 217934 36644
rect 557534 36632 557540 36644
rect 217928 36604 557540 36632
rect 217928 36592 217934 36604
rect 557534 36592 557540 36604
rect 557592 36592 557598 36644
rect 17218 36524 17224 36576
rect 17276 36564 17282 36576
rect 93946 36564 93952 36576
rect 17276 36536 93952 36564
rect 17276 36524 17282 36536
rect 93946 36524 93952 36536
rect 94004 36524 94010 36576
rect 133782 36524 133788 36576
rect 133840 36564 133846 36576
rect 164234 36564 164240 36576
rect 133840 36536 164240 36564
rect 133840 36524 133846 36536
rect 164234 36524 164240 36536
rect 164292 36524 164298 36576
rect 186222 36524 186228 36576
rect 186280 36564 186286 36576
rect 412634 36564 412640 36576
rect 186280 36536 412640 36564
rect 186280 36524 186286 36536
rect 412634 36524 412640 36536
rect 412692 36524 412698 36576
rect 422754 36524 422760 36576
rect 422812 36564 422818 36576
rect 579614 36564 579620 36576
rect 422812 36536 579620 36564
rect 422812 36524 422818 36536
rect 579614 36524 579620 36536
rect 579672 36524 579678 36576
rect 402974 35844 402980 35896
rect 403032 35884 403038 35896
rect 403342 35884 403348 35896
rect 403032 35856 403348 35884
rect 403032 35844 403038 35856
rect 403342 35844 403348 35856
rect 403400 35844 403406 35896
rect 407114 35844 407120 35896
rect 407172 35884 407178 35896
rect 408126 35884 408132 35896
rect 407172 35856 408132 35884
rect 407172 35844 407178 35856
rect 408126 35844 408132 35856
rect 408184 35844 408190 35896
rect 222378 35572 222384 35624
rect 222436 35612 222442 35624
rect 243354 35612 243360 35624
rect 222436 35584 243360 35612
rect 222436 35572 222442 35584
rect 243354 35572 243360 35584
rect 243412 35572 243418 35624
rect 251174 35572 251180 35624
rect 251232 35612 251238 35624
rect 349522 35612 349528 35624
rect 251232 35584 349528 35612
rect 251232 35572 251238 35584
rect 349522 35572 349528 35584
rect 349580 35572 349586 35624
rect 204254 35504 204260 35556
rect 204312 35544 204318 35556
rect 239398 35544 239404 35556
rect 204312 35516 239404 35544
rect 204312 35504 204318 35516
rect 239398 35504 239404 35516
rect 239456 35504 239462 35556
rect 290090 35504 290096 35556
rect 290148 35544 290154 35556
rect 434714 35544 434720 35556
rect 290148 35516 434720 35544
rect 290148 35504 290154 35516
rect 434714 35504 434720 35516
rect 434772 35504 434778 35556
rect 166994 35436 167000 35488
rect 167052 35476 167058 35488
rect 330386 35476 330392 35488
rect 167052 35448 330392 35476
rect 167052 35436 167058 35448
rect 330386 35436 330392 35448
rect 330444 35436 330450 35488
rect 171410 35368 171416 35420
rect 171468 35408 171474 35420
rect 349154 35408 349160 35420
rect 171468 35380 349160 35408
rect 171468 35368 171474 35380
rect 349154 35368 349160 35380
rect 349212 35368 349218 35420
rect 419718 35368 419724 35420
rect 419776 35408 419782 35420
rect 571334 35408 571340 35420
rect 419776 35380 571340 35408
rect 419776 35368 419782 35380
rect 571334 35368 571340 35380
rect 571392 35368 571398 35420
rect 127066 35300 127072 35352
rect 127124 35340 127130 35352
rect 222194 35340 222200 35352
rect 127124 35312 222200 35340
rect 127124 35300 127130 35312
rect 222194 35300 222200 35312
rect 222252 35300 222258 35352
rect 261202 35300 261208 35352
rect 261260 35340 261266 35352
rect 303614 35340 303620 35352
rect 261260 35312 303620 35340
rect 261260 35300 261266 35312
rect 303614 35300 303620 35312
rect 303672 35300 303678 35352
rect 311986 35300 311992 35352
rect 312044 35340 312050 35352
rect 534074 35340 534080 35352
rect 312044 35312 534080 35340
rect 312044 35300 312050 35312
rect 534074 35300 534080 35312
rect 534132 35300 534138 35352
rect 201494 35232 201500 35284
rect 201552 35272 201558 35284
rect 483014 35272 483020 35284
rect 201552 35244 483020 35272
rect 201552 35232 201558 35244
rect 483014 35232 483020 35244
rect 483072 35232 483078 35284
rect 6914 35164 6920 35216
rect 6972 35204 6978 35216
rect 41322 35204 41328 35216
rect 6972 35176 41328 35204
rect 6972 35164 6978 35176
rect 41322 35164 41328 35176
rect 41380 35164 41386 35216
rect 68922 35164 68928 35216
rect 68980 35204 68986 35216
rect 121546 35204 121552 35216
rect 68980 35176 121552 35204
rect 68980 35164 68986 35176
rect 121546 35164 121552 35176
rect 121604 35164 121610 35216
rect 219526 35164 219532 35216
rect 219584 35204 219590 35216
rect 564434 35204 564440 35216
rect 219584 35176 564440 35204
rect 219584 35164 219590 35176
rect 564434 35164 564440 35176
rect 564492 35164 564498 35216
rect 307018 34212 307024 34264
rect 307076 34252 307082 34264
rect 360378 34252 360384 34264
rect 307076 34224 360384 34252
rect 307076 34212 307082 34224
rect 360378 34212 360384 34224
rect 360436 34212 360442 34264
rect 161474 34144 161480 34196
rect 161532 34184 161538 34196
rect 230014 34184 230020 34196
rect 161532 34156 230020 34184
rect 161532 34144 161538 34156
rect 230014 34144 230020 34156
rect 230072 34144 230078 34196
rect 259454 34144 259460 34196
rect 259512 34184 259518 34196
rect 350994 34184 351000 34196
rect 259512 34156 351000 34184
rect 259512 34144 259518 34156
rect 350994 34144 351000 34156
rect 351052 34144 351058 34196
rect 140866 34076 140872 34128
rect 140924 34116 140930 34128
rect 225322 34116 225328 34128
rect 140924 34088 225328 34116
rect 140924 34076 140930 34088
rect 225322 34076 225328 34088
rect 225380 34076 225386 34128
rect 278314 34076 278320 34128
rect 278372 34116 278378 34128
rect 378226 34116 378232 34128
rect 278372 34088 378232 34116
rect 278372 34076 278378 34088
rect 378226 34076 378232 34088
rect 378284 34076 378290 34128
rect 209866 34008 209872 34060
rect 209924 34048 209930 34060
rect 340046 34048 340052 34060
rect 209924 34020 340052 34048
rect 209924 34008 209930 34020
rect 340046 34008 340052 34020
rect 340104 34008 340110 34060
rect 163682 33940 163688 33992
rect 163740 33980 163746 33992
rect 313274 33980 313280 33992
rect 163740 33952 313280 33980
rect 163740 33940 163746 33952
rect 313274 33940 313280 33952
rect 313332 33940 313338 33992
rect 408770 33940 408776 33992
rect 408828 33980 408834 33992
rect 521654 33980 521660 33992
rect 408828 33952 521660 33980
rect 408828 33940 408834 33952
rect 521654 33940 521660 33952
rect 521712 33940 521718 33992
rect 196066 33872 196072 33924
rect 196124 33912 196130 33924
rect 458174 33912 458180 33924
rect 196124 33884 458180 33912
rect 196124 33872 196130 33884
rect 458174 33872 458180 33884
rect 458232 33872 458238 33924
rect 224126 33804 224132 33856
rect 224184 33844 224190 33856
rect 489914 33844 489920 33856
rect 224184 33816 489920 33844
rect 224184 33804 224190 33816
rect 489914 33804 489920 33816
rect 489972 33804 489978 33856
rect 11054 33736 11060 33788
rect 11112 33776 11118 33788
rect 42886 33776 42892 33788
rect 11112 33748 42892 33776
rect 11112 33736 11118 33748
rect 42886 33736 42892 33748
rect 42944 33736 42950 33788
rect 55214 33736 55220 33788
rect 55272 33776 55278 33788
rect 75914 33776 75920 33788
rect 55272 33748 75920 33776
rect 55272 33736 55278 33748
rect 75914 33736 75920 33748
rect 75972 33736 75978 33788
rect 220814 33736 220820 33788
rect 220872 33776 220878 33788
rect 572714 33776 572720 33788
rect 220872 33748 572720 33776
rect 220872 33736 220878 33748
rect 572714 33736 572720 33748
rect 572772 33736 572778 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 38102 33096 38108 33108
rect 3200 33068 38108 33096
rect 3200 33056 3206 33068
rect 38102 33056 38108 33068
rect 38160 33056 38166 33108
rect 428642 33056 428648 33108
rect 428700 33096 428706 33108
rect 579890 33096 579896 33108
rect 428700 33068 579896 33096
rect 428700 33056 428706 33068
rect 579890 33056 579896 33068
rect 579948 33056 579954 33108
rect 291838 32784 291844 32836
rect 291896 32824 291902 32836
rect 357526 32824 357532 32836
rect 291896 32796 357532 32824
rect 291896 32784 291902 32796
rect 357526 32784 357532 32796
rect 357584 32784 357590 32836
rect 150618 32716 150624 32768
rect 150676 32756 150682 32768
rect 245654 32756 245660 32768
rect 150676 32728 245660 32756
rect 150676 32716 150682 32728
rect 245654 32716 245660 32728
rect 245712 32716 245718 32768
rect 275922 32716 275928 32768
rect 275980 32756 275986 32768
rect 367186 32756 367192 32768
rect 275980 32728 367192 32756
rect 275980 32716 275986 32728
rect 367186 32716 367192 32728
rect 367244 32716 367250 32768
rect 234614 32648 234620 32700
rect 234672 32688 234678 32700
rect 345014 32688 345020 32700
rect 234672 32660 345020 32688
rect 234672 32648 234678 32660
rect 345014 32648 345020 32660
rect 345072 32648 345078 32700
rect 160186 32580 160192 32632
rect 160244 32620 160250 32632
rect 295334 32620 295340 32632
rect 160244 32592 295340 32620
rect 160244 32580 160250 32592
rect 295334 32580 295340 32592
rect 295392 32580 295398 32632
rect 295978 32580 295984 32632
rect 296036 32620 296042 32632
rect 445754 32620 445760 32632
rect 296036 32592 445760 32620
rect 296036 32580 296042 32592
rect 445754 32580 445760 32592
rect 445812 32580 445818 32632
rect 181622 32512 181628 32564
rect 181680 32552 181686 32564
rect 394786 32552 394792 32564
rect 181680 32524 394792 32552
rect 181680 32512 181686 32524
rect 394786 32512 394792 32524
rect 394844 32512 394850 32564
rect 197446 32444 197452 32496
rect 197504 32484 197510 32496
rect 465166 32484 465172 32496
rect 197504 32456 465172 32484
rect 197504 32444 197510 32456
rect 465166 32444 465172 32456
rect 465224 32444 465230 32496
rect 35894 32376 35900 32428
rect 35952 32416 35958 32428
rect 47394 32416 47400 32428
rect 35952 32388 47400 32416
rect 35952 32376 35958 32388
rect 47394 32376 47400 32388
rect 47452 32376 47458 32428
rect 49878 32376 49884 32428
rect 49936 32416 49942 32428
rect 100846 32416 100852 32428
rect 49936 32388 100852 32416
rect 49936 32376 49942 32388
rect 100846 32376 100852 32388
rect 100904 32376 100910 32428
rect 216766 32376 216772 32428
rect 216824 32416 216830 32428
rect 554774 32416 554780 32428
rect 216824 32388 554780 32416
rect 216824 32376 216830 32388
rect 554774 32376 554780 32388
rect 554832 32376 554838 32428
rect 143626 31424 143632 31476
rect 143684 31464 143690 31476
rect 226334 31464 226340 31476
rect 143684 31436 226340 31464
rect 143684 31424 143690 31436
rect 226334 31424 226340 31436
rect 226392 31424 226398 31476
rect 273254 31424 273260 31476
rect 273312 31464 273318 31476
rect 353846 31464 353852 31476
rect 273312 31436 353852 31464
rect 273312 31424 273318 31436
rect 353846 31424 353852 31436
rect 353904 31424 353910 31476
rect 216674 31356 216680 31408
rect 216732 31396 216738 31408
rect 340966 31396 340972 31408
rect 216732 31368 340972 31396
rect 216732 31356 216738 31368
rect 340966 31356 340972 31368
rect 341024 31356 341030 31408
rect 133874 31288 133880 31340
rect 133932 31328 133938 31340
rect 223850 31328 223856 31340
rect 133932 31300 223856 31328
rect 133932 31288 133938 31300
rect 223850 31288 223856 31300
rect 223908 31288 223914 31340
rect 291746 31288 291752 31340
rect 291804 31328 291810 31340
rect 441614 31328 441620 31340
rect 291804 31300 441620 31328
rect 291804 31288 291810 31300
rect 441614 31288 441620 31300
rect 441672 31288 441678 31340
rect 172698 31220 172704 31272
rect 172756 31260 172762 31272
rect 345014 31260 345020 31272
rect 172756 31232 345020 31260
rect 172756 31220 172762 31232
rect 345014 31220 345020 31232
rect 345072 31220 345078 31272
rect 418246 31220 418252 31272
rect 418304 31260 418310 31272
rect 564526 31260 564532 31272
rect 418304 31232 564532 31260
rect 418304 31220 418310 31232
rect 564526 31220 564532 31232
rect 564584 31220 564590 31272
rect 20714 31152 20720 31204
rect 20772 31192 20778 31204
rect 44266 31192 44272 31204
rect 20772 31164 44272 31192
rect 20772 31152 20778 31164
rect 44266 31152 44272 31164
rect 44324 31152 44330 31204
rect 76006 31152 76012 31204
rect 76064 31152 76070 31204
rect 199562 31152 199568 31204
rect 199620 31192 199626 31204
rect 476114 31192 476120 31204
rect 199620 31164 476120 31192
rect 199620 31152 199626 31164
rect 476114 31152 476120 31164
rect 476172 31152 476178 31204
rect 44266 31016 44272 31068
rect 44324 31056 44330 31068
rect 74626 31056 74632 31068
rect 44324 31028 74632 31056
rect 44324 31016 44330 31028
rect 74626 31016 74632 31028
rect 74684 31016 74690 31068
rect 76024 31000 76052 31152
rect 206922 31084 206928 31136
rect 206980 31124 206986 31136
rect 494054 31124 494060 31136
rect 206980 31096 494060 31124
rect 206980 31084 206986 31096
rect 494054 31084 494060 31096
rect 494112 31084 494118 31136
rect 222654 31016 222660 31068
rect 222712 31056 222718 31068
rect 575474 31056 575480 31068
rect 222712 31028 575480 31056
rect 222712 31016 222718 31028
rect 575474 31016 575480 31028
rect 575532 31016 575538 31068
rect 76006 30948 76012 31000
rect 76064 30948 76070 31000
rect 276106 29996 276112 30048
rect 276164 30036 276170 30048
rect 371418 30036 371424 30048
rect 276164 30008 371424 30036
rect 276164 29996 276170 30008
rect 371418 29996 371424 30008
rect 371476 29996 371482 30048
rect 158714 29928 158720 29980
rect 158772 29968 158778 29980
rect 229094 29968 229100 29980
rect 158772 29940 229100 29968
rect 158772 29928 158778 29940
rect 229094 29928 229100 29940
rect 229152 29928 229158 29980
rect 244366 29928 244372 29980
rect 244424 29968 244430 29980
rect 347866 29968 347872 29980
rect 244424 29940 347872 29968
rect 244424 29928 244430 29940
rect 347866 29928 347872 29940
rect 347924 29928 347930 29980
rect 205634 29860 205640 29912
rect 205692 29900 205698 29912
rect 339494 29900 339500 29912
rect 205692 29872 339500 29900
rect 205692 29860 205698 29872
rect 339494 29860 339500 29872
rect 339552 29860 339558 29912
rect 405734 29860 405740 29912
rect 405792 29900 405798 29912
rect 506474 29900 506480 29912
rect 405792 29872 506480 29900
rect 405792 29860 405798 29872
rect 506474 29860 506480 29872
rect 506532 29860 506538 29912
rect 168374 29792 168380 29844
rect 168432 29832 168438 29844
rect 334158 29832 334164 29844
rect 168432 29804 334164 29832
rect 168432 29792 168438 29804
rect 334158 29792 334164 29804
rect 334216 29792 334222 29844
rect 417418 29792 417424 29844
rect 417476 29832 417482 29844
rect 560294 29832 560300 29844
rect 417476 29804 560300 29832
rect 417476 29792 417482 29804
rect 560294 29792 560300 29804
rect 560352 29792 560358 29844
rect 154758 29724 154764 29776
rect 154816 29764 154822 29776
rect 270494 29764 270500 29776
rect 154816 29736 270500 29764
rect 154816 29724 154822 29736
rect 270494 29724 270500 29736
rect 270552 29724 270558 29776
rect 309594 29724 309600 29776
rect 309652 29764 309658 29776
rect 523034 29764 523040 29776
rect 309652 29736 523040 29764
rect 309652 29724 309658 29736
rect 523034 29724 523040 29736
rect 523092 29724 523098 29776
rect 33134 29656 33140 29708
rect 33192 29696 33198 29708
rect 46934 29696 46940 29708
rect 33192 29668 46940 29696
rect 33192 29656 33198 29668
rect 46934 29656 46940 29668
rect 46992 29656 46998 29708
rect 190638 29656 190644 29708
rect 190696 29696 190702 29708
rect 426434 29696 426440 29708
rect 190696 29668 426440 29696
rect 190696 29656 190702 29668
rect 426434 29656 426440 29668
rect 426492 29656 426498 29708
rect 15838 29588 15844 29640
rect 15896 29628 15902 29640
rect 92658 29628 92664 29640
rect 15896 29600 92664 29628
rect 15896 29588 15902 29600
rect 92658 29588 92664 29600
rect 92716 29588 92722 29640
rect 205082 29588 205088 29640
rect 205140 29628 205146 29640
rect 500954 29628 500960 29640
rect 205140 29600 500960 29628
rect 205140 29588 205146 29600
rect 500954 29588 500960 29600
rect 501012 29588 501018 29640
rect 262766 28704 262772 28756
rect 262824 28744 262830 28756
rect 310514 28744 310520 28756
rect 262824 28716 310520 28744
rect 262824 28704 262830 28716
rect 310514 28704 310520 28716
rect 310572 28704 310578 28756
rect 262214 28636 262220 28688
rect 262272 28676 262278 28688
rect 352006 28676 352012 28688
rect 262272 28648 352012 28676
rect 262272 28636 262278 28648
rect 352006 28636 352012 28648
rect 352064 28636 352070 28688
rect 279234 28568 279240 28620
rect 279292 28608 279298 28620
rect 385218 28608 385224 28620
rect 279292 28580 385224 28608
rect 279292 28568 279298 28580
rect 385218 28568 385224 28580
rect 385276 28568 385282 28620
rect 165706 28500 165712 28552
rect 165764 28540 165770 28552
rect 320358 28540 320364 28552
rect 165764 28512 320364 28540
rect 165764 28500 165770 28512
rect 320358 28500 320364 28512
rect 320416 28500 320422 28552
rect 176746 28432 176752 28484
rect 176804 28472 176810 28484
rect 333054 28472 333060 28484
rect 176804 28444 333060 28472
rect 176804 28432 176810 28444
rect 333054 28432 333060 28444
rect 333112 28432 333118 28484
rect 404446 28432 404452 28484
rect 404504 28472 404510 28484
rect 499574 28472 499580 28484
rect 404504 28444 499580 28472
rect 404504 28432 404510 28444
rect 499574 28432 499580 28444
rect 499632 28432 499638 28484
rect 151814 28364 151820 28416
rect 151872 28404 151878 28416
rect 259638 28404 259644 28416
rect 151872 28376 259644 28404
rect 151872 28364 151878 28376
rect 259638 28364 259644 28376
rect 259696 28364 259702 28416
rect 309778 28364 309784 28416
rect 309836 28404 309842 28416
rect 513374 28404 513380 28416
rect 309836 28376 513380 28404
rect 309836 28364 309842 28376
rect 513374 28364 513380 28376
rect 513432 28364 513438 28416
rect 183922 28296 183928 28348
rect 183980 28336 183986 28348
rect 405734 28336 405740 28348
rect 183980 28308 405740 28336
rect 183980 28296 183986 28308
rect 405734 28296 405740 28308
rect 405792 28296 405798 28348
rect 415762 28296 415768 28348
rect 415820 28336 415826 28348
rect 553394 28336 553400 28348
rect 415820 28308 553400 28336
rect 415820 28296 415826 28308
rect 553394 28296 553400 28308
rect 553452 28296 553458 28348
rect 2774 28228 2780 28280
rect 2832 28268 2838 28280
rect 66898 28268 66904 28280
rect 2832 28240 66904 28268
rect 2832 28228 2838 28240
rect 66898 28228 66904 28240
rect 66956 28228 66962 28280
rect 209038 28228 209044 28280
rect 209096 28268 209102 28280
rect 507854 28268 507860 28280
rect 209096 28240 507860 28268
rect 209096 28228 209102 28240
rect 507854 28228 507860 28240
rect 507912 28228 507918 28280
rect 293954 27344 293960 27396
rect 294012 27384 294018 27396
rect 356698 27384 356704 27396
rect 294012 27356 356704 27384
rect 294012 27344 294018 27356
rect 356698 27344 356704 27356
rect 356756 27344 356762 27396
rect 273714 27276 273720 27328
rect 273772 27316 273778 27328
rect 360194 27316 360200 27328
rect 273772 27288 360200 27316
rect 273772 27276 273778 27288
rect 360194 27276 360200 27288
rect 360252 27276 360258 27328
rect 294138 27208 294144 27260
rect 294196 27248 294202 27260
rect 452654 27248 452660 27260
rect 294196 27220 452660 27248
rect 294196 27208 294202 27220
rect 452654 27208 452660 27220
rect 452712 27208 452718 27260
rect 167546 27140 167552 27192
rect 167604 27180 167610 27192
rect 331214 27180 331220 27192
rect 167604 27152 331220 27180
rect 167604 27140 167610 27152
rect 331214 27140 331220 27152
rect 331272 27140 331278 27192
rect 140038 27072 140044 27124
rect 140096 27112 140102 27124
rect 323762 27112 323768 27124
rect 140096 27084 323768 27112
rect 140096 27072 140102 27084
rect 323762 27072 323768 27084
rect 323820 27072 323826 27124
rect 412818 27072 412824 27124
rect 412876 27112 412882 27124
rect 539594 27112 539600 27124
rect 412876 27084 539600 27112
rect 412876 27072 412882 27084
rect 539594 27072 539600 27084
rect 539652 27072 539658 27124
rect 67818 27004 67824 27056
rect 67876 27044 67882 27056
rect 104066 27044 104072 27056
rect 67876 27016 104072 27044
rect 67876 27004 67882 27016
rect 104066 27004 104072 27016
rect 104124 27004 104130 27056
rect 153562 27004 153568 27056
rect 153620 27044 153626 27056
rect 267826 27044 267832 27056
rect 153620 27016 267832 27044
rect 153620 27004 153626 27016
rect 267826 27004 267832 27016
rect 267884 27004 267890 27056
rect 309134 27004 309140 27056
rect 309192 27044 309198 27056
rect 520274 27044 520280 27056
rect 309192 27016 520280 27044
rect 309192 27004 309198 27016
rect 520274 27004 520280 27016
rect 520332 27004 520338 27056
rect 187050 26936 187056 26988
rect 187108 26976 187114 26988
rect 419534 26976 419540 26988
rect 187108 26948 419540 26976
rect 187108 26936 187114 26948
rect 419534 26936 419540 26948
rect 419592 26936 419598 26988
rect 14458 26868 14464 26920
rect 14516 26908 14522 26920
rect 67634 26908 67640 26920
rect 14516 26880 67640 26908
rect 14516 26868 14522 26880
rect 67634 26868 67640 26880
rect 67692 26868 67698 26920
rect 207382 26868 207388 26920
rect 207440 26908 207446 26920
rect 511994 26908 512000 26920
rect 207440 26880 512000 26908
rect 207440 26868 207446 26880
rect 511994 26868 512000 26880
rect 512052 26868 512058 26920
rect 151814 25916 151820 25968
rect 151872 25956 151878 25968
rect 227806 25956 227812 25968
rect 151872 25928 227812 25956
rect 151872 25916 151878 25928
rect 227806 25916 227812 25928
rect 227864 25916 227870 25968
rect 248598 25916 248604 25968
rect 248656 25956 248662 25968
rect 330570 25956 330576 25968
rect 248656 25928 330576 25956
rect 248656 25916 248662 25928
rect 330570 25916 330576 25928
rect 330628 25916 330634 25968
rect 201494 25848 201500 25900
rect 201552 25888 201558 25900
rect 338206 25888 338212 25900
rect 201552 25860 338212 25888
rect 201552 25848 201558 25860
rect 338206 25848 338212 25860
rect 338264 25848 338270 25900
rect 143718 25780 143724 25832
rect 143776 25820 143782 25832
rect 220814 25820 220820 25832
rect 143776 25792 220820 25820
rect 143776 25780 143782 25792
rect 220814 25780 220820 25792
rect 220872 25780 220878 25832
rect 294046 25780 294052 25832
rect 294104 25820 294110 25832
rect 456886 25820 456892 25832
rect 294104 25792 456892 25820
rect 294104 25780 294110 25792
rect 456886 25780 456892 25792
rect 456944 25780 456950 25832
rect 218698 25712 218704 25764
rect 218756 25752 218762 25764
rect 390646 25752 390652 25764
rect 218756 25724 390652 25752
rect 218756 25712 218762 25724
rect 390646 25712 390652 25724
rect 390704 25712 390710 25764
rect 421006 25712 421012 25764
rect 421064 25752 421070 25764
rect 574094 25752 574100 25764
rect 421064 25724 574100 25752
rect 421064 25712 421070 25724
rect 574094 25712 574100 25724
rect 574152 25712 574158 25764
rect 158806 25644 158812 25696
rect 158864 25684 158870 25696
rect 292574 25684 292580 25696
rect 158864 25656 292580 25684
rect 158864 25644 158870 25656
rect 292574 25644 292580 25656
rect 292632 25644 292638 25696
rect 314654 25644 314660 25696
rect 314712 25684 314718 25696
rect 547874 25684 547880 25696
rect 314712 25656 547880 25684
rect 314712 25644 314718 25656
rect 547874 25644 547880 25656
rect 547932 25644 547938 25696
rect 193214 25576 193220 25628
rect 193272 25616 193278 25628
rect 451274 25616 451280 25628
rect 193272 25588 451280 25616
rect 193272 25576 193278 25588
rect 451274 25576 451280 25588
rect 451332 25576 451338 25628
rect 17954 25508 17960 25560
rect 18012 25548 18018 25560
rect 69014 25548 69020 25560
rect 18012 25520 69020 25548
rect 18012 25508 18018 25520
rect 69014 25508 69020 25520
rect 69072 25508 69078 25560
rect 77294 25508 77300 25560
rect 77352 25548 77358 25560
rect 106366 25548 106372 25560
rect 77352 25520 106372 25548
rect 77352 25508 77358 25520
rect 106366 25508 106372 25520
rect 106424 25508 106430 25560
rect 214006 25508 214012 25560
rect 214064 25548 214070 25560
rect 543734 25548 543740 25560
rect 214064 25520 543740 25548
rect 214064 25508 214070 25520
rect 543734 25508 543740 25520
rect 543792 25508 543798 25560
rect 149054 24488 149060 24540
rect 149112 24528 149118 24540
rect 249978 24528 249984 24540
rect 149112 24500 249984 24528
rect 149112 24488 149118 24500
rect 249978 24488 249984 24500
rect 250036 24488 250042 24540
rect 276014 24488 276020 24540
rect 276072 24528 276078 24540
rect 353938 24528 353944 24540
rect 276072 24500 353944 24528
rect 276072 24488 276078 24500
rect 353938 24488 353944 24500
rect 353996 24488 354002 24540
rect 241606 24420 241612 24472
rect 241664 24460 241670 24472
rect 346486 24460 346492 24472
rect 241664 24432 346492 24460
rect 241664 24420 241670 24432
rect 346486 24420 346492 24432
rect 346544 24420 346550 24472
rect 184934 24352 184940 24404
rect 184992 24392 184998 24404
rect 333974 24392 333980 24404
rect 184992 24364 333980 24392
rect 184992 24352 184998 24364
rect 333974 24352 333980 24364
rect 334032 24352 334038 24404
rect 182174 24284 182180 24336
rect 182232 24324 182238 24336
rect 398926 24324 398932 24336
rect 182232 24296 398932 24324
rect 182232 24284 182238 24296
rect 398926 24284 398932 24296
rect 398984 24284 398990 24336
rect 412726 24284 412732 24336
rect 412784 24324 412790 24336
rect 542354 24324 542360 24336
rect 412784 24296 542360 24324
rect 412784 24284 412790 24296
rect 542354 24284 542360 24296
rect 542412 24284 542418 24336
rect 170398 24216 170404 24268
rect 170456 24256 170462 24268
rect 309134 24256 309140 24268
rect 170456 24228 309140 24256
rect 170456 24216 170462 24228
rect 309134 24216 309140 24228
rect 309192 24216 309198 24268
rect 318794 24216 318800 24268
rect 318852 24256 318858 24268
rect 565814 24256 565820 24268
rect 318852 24228 565820 24256
rect 318852 24216 318858 24228
rect 565814 24216 565820 24228
rect 565872 24216 565878 24268
rect 70578 24148 70584 24200
rect 70636 24188 70642 24200
rect 104894 24188 104900 24200
rect 70636 24160 104900 24188
rect 70636 24148 70642 24160
rect 104894 24148 104900 24160
rect 104952 24148 104958 24200
rect 197354 24148 197360 24200
rect 197412 24188 197418 24200
rect 469214 24188 469220 24200
rect 197412 24160 469220 24188
rect 197412 24148 197418 24160
rect 469214 24148 469220 24160
rect 469272 24148 469278 24200
rect 22094 24080 22100 24132
rect 22152 24120 22158 24132
rect 70486 24120 70492 24132
rect 22152 24092 70492 24120
rect 22152 24080 22158 24092
rect 70486 24080 70492 24092
rect 70544 24080 70550 24132
rect 209958 24080 209964 24132
rect 210016 24120 210022 24132
rect 523126 24120 523132 24132
rect 210016 24092 523132 24120
rect 210016 24080 210022 24092
rect 523126 24080 523132 24092
rect 523184 24080 523190 24132
rect 263778 23196 263784 23248
rect 263836 23236 263842 23248
rect 314654 23236 314660 23248
rect 263836 23208 314660 23236
rect 263836 23196 263842 23208
rect 314654 23196 314660 23208
rect 314712 23196 314718 23248
rect 266538 23128 266544 23180
rect 266596 23168 266602 23180
rect 351914 23168 351920 23180
rect 266596 23140 351920 23168
rect 266596 23128 266602 23140
rect 351914 23128 351920 23140
rect 351972 23128 351978 23180
rect 288526 23060 288532 23112
rect 288584 23100 288590 23112
rect 427814 23100 427820 23112
rect 288584 23072 427820 23100
rect 288584 23060 288590 23072
rect 427814 23060 427820 23072
rect 427872 23060 427878 23112
rect 194686 22992 194692 23044
rect 194744 23032 194750 23044
rect 336734 23032 336740 23044
rect 194744 23004 336740 23032
rect 194744 22992 194750 23004
rect 336734 22992 336740 23004
rect 336792 22992 336798 23044
rect 165614 22924 165620 22976
rect 165672 22964 165678 22976
rect 324314 22964 324320 22976
rect 165672 22936 324320 22964
rect 165672 22924 165678 22936
rect 324314 22924 324320 22936
rect 324372 22924 324378 22976
rect 407206 22924 407212 22976
rect 407264 22964 407270 22976
rect 514754 22964 514760 22976
rect 407264 22936 514760 22964
rect 407264 22924 407270 22936
rect 514754 22924 514760 22936
rect 514812 22924 514818 22976
rect 151906 22856 151912 22908
rect 151964 22896 151970 22908
rect 263686 22896 263692 22908
rect 151964 22868 263692 22896
rect 151964 22856 151970 22868
rect 263686 22856 263692 22868
rect 263744 22856 263750 22908
rect 307754 22856 307760 22908
rect 307812 22896 307818 22908
rect 516134 22896 516140 22908
rect 307812 22868 516140 22896
rect 307812 22856 307818 22868
rect 516134 22856 516140 22868
rect 516192 22856 516198 22908
rect 34514 22788 34520 22840
rect 34572 22828 34578 22840
rect 71866 22828 71872 22840
rect 34572 22800 71872 22828
rect 34572 22788 34578 22800
rect 71866 22788 71872 22800
rect 71924 22788 71930 22840
rect 188338 22788 188344 22840
rect 188396 22828 188402 22840
rect 408494 22828 408500 22840
rect 188396 22800 408500 22828
rect 188396 22788 188402 22800
rect 408494 22788 408500 22800
rect 408552 22788 408558 22840
rect 418154 22788 418160 22840
rect 418212 22828 418218 22840
rect 567194 22828 567200 22840
rect 418212 22800 567200 22828
rect 418212 22788 418218 22800
rect 567194 22788 567200 22800
rect 567252 22788 567258 22840
rect 63586 22720 63592 22772
rect 63644 22760 63650 22772
rect 103514 22760 103520 22772
rect 63644 22732 103520 22760
rect 63644 22720 63650 22732
rect 103514 22720 103520 22732
rect 103572 22720 103578 22772
rect 205726 22720 205732 22772
rect 205784 22760 205790 22772
rect 505094 22760 505100 22772
rect 205784 22732 505100 22760
rect 205784 22720 205790 22732
rect 505094 22720 505100 22732
rect 505152 22720 505158 22772
rect 294598 21836 294604 21888
rect 294656 21876 294662 21888
rect 357434 21876 357440 21888
rect 294656 21848 357440 21876
rect 294656 21836 294662 21848
rect 357434 21836 357440 21848
rect 357492 21836 357498 21888
rect 280798 21768 280804 21820
rect 280856 21808 280862 21820
rect 382366 21808 382372 21820
rect 280856 21780 382372 21808
rect 280856 21768 280862 21780
rect 382366 21768 382372 21780
rect 382424 21768 382430 21820
rect 219526 21700 219532 21752
rect 219584 21740 219590 21752
rect 342254 21740 342260 21752
rect 219584 21712 342260 21740
rect 219584 21700 219590 21712
rect 342254 21700 342260 21712
rect 342312 21700 342318 21752
rect 262306 21632 262312 21684
rect 262364 21672 262370 21684
rect 307754 21672 307760 21684
rect 262364 21644 307760 21672
rect 262364 21632 262370 21644
rect 307754 21632 307760 21644
rect 307812 21632 307818 21684
rect 312538 21632 312544 21684
rect 312596 21672 312602 21684
rect 463694 21672 463700 21684
rect 312596 21644 463700 21672
rect 312596 21632 312602 21644
rect 463694 21632 463700 21644
rect 463752 21632 463758 21684
rect 164326 21564 164332 21616
rect 164384 21604 164390 21616
rect 316218 21604 316224 21616
rect 164384 21576 316224 21604
rect 164384 21564 164390 21576
rect 316218 21564 316224 21576
rect 316276 21564 316282 21616
rect 150526 21496 150532 21548
rect 150584 21536 150590 21548
rect 256878 21536 256884 21548
rect 150584 21508 256884 21536
rect 150584 21496 150590 21508
rect 256878 21496 256884 21508
rect 256936 21496 256942 21548
rect 306374 21496 306380 21548
rect 306432 21536 306438 21548
rect 509234 21536 509240 21548
rect 306432 21508 509240 21536
rect 306432 21496 306438 21508
rect 509234 21496 509240 21508
rect 509292 21496 509298 21548
rect 27614 21428 27620 21480
rect 27672 21468 27678 21480
rect 70394 21468 70400 21480
rect 27672 21440 70400 21468
rect 27672 21428 27678 21440
rect 70394 21428 70400 21440
rect 70452 21428 70458 21480
rect 183554 21428 183560 21480
rect 183612 21468 183618 21480
rect 401686 21468 401692 21480
rect 183612 21440 401692 21468
rect 183612 21428 183618 21440
rect 401686 21428 401692 21440
rect 401744 21428 401750 21480
rect 409966 21428 409972 21480
rect 410024 21468 410030 21480
rect 528554 21468 528560 21480
rect 410024 21440 528560 21468
rect 410024 21428 410030 21440
rect 528554 21428 528560 21440
rect 528612 21428 528618 21480
rect 56778 21360 56784 21412
rect 56836 21400 56842 21412
rect 101398 21400 101404 21412
rect 56836 21372 101404 21400
rect 56836 21360 56842 21372
rect 101398 21360 101404 21372
rect 101456 21360 101462 21412
rect 129734 21360 129740 21412
rect 129792 21400 129798 21412
rect 157334 21400 157340 21412
rect 129792 21372 157340 21400
rect 129792 21360 129798 21372
rect 157334 21360 157340 21372
rect 157392 21360 157398 21412
rect 204346 21360 204352 21412
rect 204404 21400 204410 21412
rect 498194 21400 498200 21412
rect 204404 21372 498200 21400
rect 204404 21360 204410 21372
rect 498194 21360 498200 21372
rect 498252 21360 498258 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 38010 20652 38016 20664
rect 3476 20624 38016 20652
rect 3476 20612 3482 20624
rect 38010 20612 38016 20624
rect 38068 20612 38074 20664
rect 428550 20612 428556 20664
rect 428608 20652 428614 20664
rect 579890 20652 579896 20664
rect 428608 20624 579896 20652
rect 428608 20612 428614 20624
rect 579890 20612 579896 20624
rect 579948 20612 579954 20664
rect 267918 20340 267924 20392
rect 267976 20380 267982 20392
rect 332594 20380 332600 20392
rect 267976 20352 332600 20380
rect 267976 20340 267982 20352
rect 332594 20340 332600 20352
rect 332652 20340 332658 20392
rect 307110 20272 307116 20324
rect 307168 20312 307174 20324
rect 374178 20312 374184 20324
rect 307168 20284 374184 20312
rect 307168 20272 307174 20284
rect 374178 20272 374184 20284
rect 374236 20272 374242 20324
rect 237558 20204 237564 20256
rect 237616 20244 237622 20256
rect 346394 20244 346400 20256
rect 237616 20216 346400 20244
rect 237616 20204 237622 20216
rect 346394 20204 346400 20216
rect 346452 20204 346458 20256
rect 200758 20136 200764 20188
rect 200816 20176 200822 20188
rect 338206 20176 338212 20188
rect 200816 20148 338212 20176
rect 200816 20136 200822 20148
rect 338206 20136 338212 20148
rect 338264 20136 338270 20188
rect 409874 20136 409880 20188
rect 409932 20176 409938 20188
rect 524414 20176 524420 20188
rect 409932 20148 524420 20176
rect 409932 20136 409938 20148
rect 524414 20136 524420 20148
rect 524472 20136 524478 20188
rect 157518 20068 157524 20120
rect 157576 20108 157582 20120
rect 284478 20108 284484 20120
rect 157576 20080 284484 20108
rect 157576 20068 157582 20080
rect 284478 20068 284484 20080
rect 284536 20068 284542 20120
rect 288434 20068 288440 20120
rect 288492 20108 288498 20120
rect 432046 20108 432052 20120
rect 288492 20080 432052 20108
rect 288492 20068 288498 20080
rect 432046 20068 432052 20080
rect 432104 20068 432110 20120
rect 52638 20000 52644 20052
rect 52696 20040 52702 20052
rect 76006 20040 76012 20052
rect 52696 20012 76012 20040
rect 52696 20000 52702 20012
rect 76006 20000 76012 20012
rect 76064 20000 76070 20052
rect 189074 20000 189080 20052
rect 189132 20040 189138 20052
rect 430574 20040 430580 20052
rect 189132 20012 430580 20040
rect 189132 20000 189138 20012
rect 430574 20000 430580 20012
rect 430632 20000 430638 20052
rect 74626 19932 74632 19984
rect 74684 19972 74690 19984
rect 104158 19972 104164 19984
rect 74684 19944 104164 19972
rect 74684 19932 74690 19944
rect 104158 19932 104164 19944
rect 104216 19932 104222 19984
rect 139486 19932 139492 19984
rect 139544 19972 139550 19984
rect 207014 19972 207020 19984
rect 139544 19944 207020 19972
rect 139544 19932 139550 19944
rect 207014 19932 207020 19944
rect 207072 19932 207078 19984
rect 215294 19932 215300 19984
rect 215352 19972 215358 19984
rect 550634 19972 550640 19984
rect 215352 19944 550640 19972
rect 215352 19932 215358 19944
rect 550634 19932 550640 19944
rect 550692 19932 550698 19984
rect 255498 18980 255504 19032
rect 255556 19020 255562 19032
rect 348418 19020 348424 19032
rect 255556 18992 348424 19020
rect 255556 18980 255562 18992
rect 348418 18980 348424 18992
rect 348476 18980 348482 19032
rect 139394 18912 139400 18964
rect 139452 18952 139458 18964
rect 202874 18952 202880 18964
rect 139452 18924 202880 18952
rect 139452 18912 139458 18924
rect 202874 18912 202880 18924
rect 202932 18912 202938 18964
rect 280246 18912 280252 18964
rect 280304 18952 280310 18964
rect 389358 18952 389364 18964
rect 280304 18924 389364 18952
rect 280304 18912 280310 18924
rect 389358 18912 389364 18924
rect 389416 18912 389422 18964
rect 174078 18844 174084 18896
rect 174136 18884 174142 18896
rect 330478 18884 330484 18896
rect 174136 18856 330484 18884
rect 174136 18844 174142 18856
rect 330478 18844 330484 18856
rect 330536 18844 330542 18896
rect 172606 18776 172612 18828
rect 172664 18816 172670 18828
rect 351914 18816 351920 18828
rect 172664 18788 351920 18816
rect 172664 18776 172670 18788
rect 351914 18776 351920 18788
rect 351972 18776 351978 18828
rect 407114 18776 407120 18828
rect 407172 18816 407178 18828
rect 517514 18816 517520 18828
rect 407172 18788 517520 18816
rect 407172 18776 407178 18788
rect 517514 18776 517520 18788
rect 517572 18776 517578 18828
rect 157426 18708 157432 18760
rect 157484 18748 157490 18760
rect 288434 18748 288440 18760
rect 157484 18720 288440 18748
rect 157484 18708 157490 18720
rect 288434 18708 288440 18720
rect 288492 18708 288498 18760
rect 310606 18708 310612 18760
rect 310664 18748 310670 18760
rect 527174 18748 527180 18760
rect 310664 18720 527180 18748
rect 310664 18708 310670 18720
rect 527174 18708 527180 18720
rect 527232 18708 527238 18760
rect 48314 18640 48320 18692
rect 48372 18680 48378 18692
rect 74534 18680 74540 18692
rect 48372 18652 74540 18680
rect 48372 18640 48378 18652
rect 74534 18640 74540 18652
rect 74592 18640 74598 18692
rect 195238 18640 195244 18692
rect 195296 18680 195302 18692
rect 448514 18680 448520 18692
rect 195296 18652 448520 18680
rect 195296 18640 195302 18652
rect 448514 18640 448520 18652
rect 448572 18640 448578 18692
rect 60918 18572 60924 18624
rect 60976 18612 60982 18624
rect 102226 18612 102232 18624
rect 60976 18584 102232 18612
rect 60976 18572 60982 18584
rect 102226 18572 102232 18584
rect 102284 18572 102290 18624
rect 201586 18572 201592 18624
rect 201644 18612 201650 18624
rect 487154 18612 487160 18624
rect 201644 18584 487160 18612
rect 201644 18572 201650 18584
rect 487154 18572 487160 18584
rect 487212 18572 487218 18624
rect 269298 17620 269304 17672
rect 269356 17660 269362 17672
rect 353294 17660 353300 17672
rect 269356 17632 353300 17660
rect 269356 17620 269362 17632
rect 353294 17620 353300 17632
rect 353352 17620 353358 17672
rect 212718 17552 212724 17604
rect 212776 17592 212782 17604
rect 340138 17592 340144 17604
rect 212776 17564 340144 17592
rect 212776 17552 212782 17564
rect 340138 17552 340144 17564
rect 340196 17552 340202 17604
rect 136818 17484 136824 17536
rect 136876 17524 136882 17536
rect 224218 17524 224224 17536
rect 136876 17496 224224 17524
rect 136876 17484 136882 17496
rect 224218 17484 224224 17496
rect 224276 17484 224282 17536
rect 291194 17484 291200 17536
rect 291252 17524 291258 17536
rect 438854 17524 438860 17536
rect 291252 17496 438860 17524
rect 291252 17484 291258 17496
rect 438854 17484 438860 17496
rect 438912 17484 438918 17536
rect 169754 17416 169760 17468
rect 169812 17456 169818 17468
rect 340966 17456 340972 17468
rect 169812 17428 340972 17456
rect 169812 17416 169818 17428
rect 340966 17416 340972 17428
rect 341024 17416 341030 17468
rect 416774 17416 416780 17468
rect 416832 17456 416838 17468
rect 556154 17456 556160 17468
rect 416832 17428 556160 17456
rect 416832 17416 416838 17428
rect 556154 17416 556160 17428
rect 556212 17416 556218 17468
rect 195974 17348 195980 17400
rect 196032 17388 196038 17400
rect 462314 17388 462320 17400
rect 196032 17360 462320 17388
rect 196032 17348 196038 17360
rect 462314 17348 462320 17360
rect 462372 17348 462378 17400
rect 66254 17280 66260 17332
rect 66312 17320 66318 17332
rect 78766 17320 78772 17332
rect 66312 17292 78772 17320
rect 66312 17280 66318 17292
rect 78766 17280 78772 17292
rect 78824 17280 78830 17332
rect 200114 17280 200120 17332
rect 200172 17320 200178 17332
rect 480254 17320 480260 17332
rect 200172 17292 480260 17320
rect 200172 17280 200178 17292
rect 480254 17280 480260 17292
rect 480312 17280 480318 17332
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 67726 17252 67732 17264
rect 8352 17224 67732 17252
rect 8352 17212 8358 17224
rect 67726 17212 67732 17224
rect 67784 17212 67790 17264
rect 88426 17212 88432 17264
rect 88484 17252 88490 17264
rect 104894 17252 104900 17264
rect 88484 17224 104900 17252
rect 88484 17212 88490 17224
rect 104894 17212 104900 17224
rect 104952 17212 104958 17264
rect 134058 17212 134064 17264
rect 134116 17252 134122 17264
rect 182174 17252 182180 17264
rect 134116 17224 182180 17252
rect 134116 17212 134122 17224
rect 182174 17212 182180 17224
rect 182232 17212 182238 17264
rect 219434 17212 219440 17264
rect 219492 17252 219498 17264
rect 568574 17252 568580 17264
rect 219492 17224 568580 17252
rect 219492 17212 219498 17224
rect 568574 17212 568580 17224
rect 568632 17212 568638 17264
rect 298278 16396 298284 16448
rect 298336 16436 298342 16448
rect 358906 16436 358912 16448
rect 298336 16408 358912 16436
rect 298336 16396 298342 16408
rect 358906 16396 358912 16408
rect 358964 16396 358970 16448
rect 227530 16328 227536 16380
rect 227588 16368 227594 16380
rect 343726 16368 343732 16380
rect 227588 16340 343732 16368
rect 227588 16328 227594 16340
rect 343726 16328 343732 16340
rect 343784 16328 343790 16380
rect 198734 16260 198740 16312
rect 198792 16300 198798 16312
rect 338114 16300 338120 16312
rect 198792 16272 338120 16300
rect 198792 16260 198798 16272
rect 338114 16260 338120 16272
rect 338172 16260 338178 16312
rect 331858 16192 331864 16244
rect 331916 16232 331922 16244
rect 473446 16232 473452 16244
rect 331916 16204 473452 16232
rect 331916 16192 331922 16204
rect 473446 16192 473452 16204
rect 473504 16192 473510 16244
rect 192018 16124 192024 16176
rect 192076 16164 192082 16176
rect 335354 16164 335360 16176
rect 192076 16136 335360 16164
rect 192076 16124 192082 16136
rect 335354 16124 335360 16136
rect 335412 16124 335418 16176
rect 188522 16056 188528 16108
rect 188580 16096 188586 16108
rect 335446 16096 335452 16108
rect 188580 16068 335452 16096
rect 188580 16056 188586 16068
rect 335446 16056 335452 16068
rect 335504 16056 335510 16108
rect 292666 15988 292672 16040
rect 292724 16028 292730 16040
rect 448606 16028 448612 16040
rect 292724 16000 448612 16028
rect 292724 15988 292730 16000
rect 448606 15988 448612 16000
rect 448664 15988 448670 16040
rect 81618 15920 81624 15972
rect 81676 15960 81682 15972
rect 107746 15960 107752 15972
rect 81676 15932 107752 15960
rect 81676 15920 81682 15932
rect 107746 15920 107752 15932
rect 107804 15920 107810 15972
rect 133966 15920 133972 15972
rect 134024 15960 134030 15972
rect 178586 15960 178592 15972
rect 134024 15932 178592 15960
rect 134024 15920 134030 15932
rect 178586 15920 178592 15932
rect 178644 15920 178650 15972
rect 180978 15920 180984 15972
rect 181036 15960 181042 15972
rect 334066 15960 334072 15972
rect 181036 15932 334072 15960
rect 181036 15920 181042 15932
rect 334066 15920 334072 15932
rect 334124 15920 334130 15972
rect 342898 15920 342904 15972
rect 342956 15960 342962 15972
rect 547966 15960 547972 15972
rect 342956 15932 547972 15960
rect 342956 15920 342962 15932
rect 547966 15920 547972 15932
rect 548024 15920 548030 15972
rect 59354 15852 59360 15904
rect 59412 15892 59418 15904
rect 93946 15892 93952 15904
rect 59412 15864 93952 15892
rect 59412 15852 59418 15864
rect 93946 15852 93952 15864
rect 94004 15852 94010 15904
rect 147858 15852 147864 15904
rect 147916 15892 147922 15904
rect 226426 15892 226432 15904
rect 147916 15864 226432 15892
rect 147916 15852 147922 15864
rect 226426 15852 226432 15864
rect 226484 15852 226490 15904
rect 318058 15852 318064 15904
rect 318116 15892 318122 15904
rect 545482 15892 545488 15904
rect 318116 15864 545488 15892
rect 318116 15852 318122 15864
rect 545482 15852 545488 15864
rect 545540 15852 545546 15904
rect 262858 14968 262864 15020
rect 262916 15008 262922 15020
rect 300762 15008 300768 15020
rect 262916 14980 300768 15008
rect 262916 14968 262922 14980
rect 300762 14968 300768 14980
rect 300820 14968 300826 15020
rect 280706 14900 280712 14952
rect 280764 14940 280770 14952
rect 356146 14940 356152 14952
rect 280764 14912 356152 14940
rect 280764 14900 280770 14912
rect 356146 14900 356152 14912
rect 356204 14900 356210 14952
rect 231026 14832 231032 14884
rect 231084 14872 231090 14884
rect 345106 14872 345112 14884
rect 231084 14844 345112 14872
rect 231084 14832 231090 14844
rect 345106 14832 345112 14844
rect 345164 14832 345170 14884
rect 170306 14764 170312 14816
rect 170364 14804 170370 14816
rect 331306 14804 331312 14816
rect 170364 14776 331312 14804
rect 170364 14764 170370 14776
rect 331306 14764 331312 14776
rect 331364 14764 331370 14816
rect 218054 14696 218060 14748
rect 218112 14736 218118 14748
rect 242158 14736 242164 14748
rect 218112 14708 242164 14736
rect 218112 14696 218118 14708
rect 242158 14696 242164 14708
rect 242216 14696 242222 14748
rect 295426 14696 295432 14748
rect 295484 14736 295490 14748
rect 459922 14736 459928 14748
rect 295484 14708 459928 14736
rect 295484 14696 295490 14708
rect 459922 14696 459928 14708
rect 459980 14696 459986 14748
rect 211706 14628 211712 14680
rect 211764 14668 211770 14680
rect 240226 14668 240232 14680
rect 211764 14640 240232 14668
rect 211764 14628 211770 14640
rect 240226 14628 240232 14640
rect 240284 14628 240290 14680
rect 298186 14628 298192 14680
rect 298244 14668 298250 14680
rect 470594 14668 470600 14680
rect 298244 14640 470600 14668
rect 298244 14628 298250 14640
rect 470594 14628 470600 14640
rect 470652 14628 470658 14680
rect 193214 14560 193220 14612
rect 193272 14600 193278 14612
rect 237466 14600 237472 14612
rect 193272 14572 237472 14600
rect 193272 14560 193278 14572
rect 237466 14560 237472 14572
rect 237524 14560 237530 14612
rect 298094 14560 298100 14612
rect 298152 14600 298158 14612
rect 474090 14600 474096 14612
rect 298152 14572 474096 14600
rect 298152 14560 298158 14572
rect 474090 14560 474096 14572
rect 474148 14560 474154 14612
rect 30834 14492 30840 14544
rect 30892 14532 30898 14544
rect 71774 14532 71780 14544
rect 30892 14504 71780 14532
rect 30892 14492 30898 14504
rect 71774 14492 71780 14504
rect 71832 14492 71838 14544
rect 128998 14492 129004 14544
rect 129056 14532 129062 14544
rect 150618 14532 150624 14544
rect 129056 14504 150624 14532
rect 129056 14492 129062 14504
rect 150618 14492 150624 14504
rect 150676 14492 150682 14544
rect 155954 14492 155960 14544
rect 156012 14532 156018 14544
rect 281718 14532 281724 14544
rect 156012 14504 281724 14532
rect 156012 14492 156018 14504
rect 281718 14492 281724 14504
rect 281776 14492 281782 14544
rect 299566 14492 299572 14544
rect 299624 14532 299630 14544
rect 478138 14532 478144 14544
rect 299624 14504 478144 14532
rect 299624 14492 299630 14504
rect 478138 14492 478144 14504
rect 478196 14492 478202 14544
rect 64966 14424 64972 14476
rect 65024 14464 65030 14476
rect 114738 14464 114744 14476
rect 65024 14436 114744 14464
rect 65024 14424 65030 14436
rect 114738 14424 114744 14436
rect 114796 14424 114802 14476
rect 129090 14424 129096 14476
rect 129148 14464 129154 14476
rect 321554 14464 321560 14476
rect 129148 14436 321560 14464
rect 129148 14424 129154 14436
rect 321554 14424 321560 14436
rect 321612 14424 321618 14476
rect 414014 14424 414020 14476
rect 414072 14464 414078 14476
rect 546494 14464 546500 14476
rect 414072 14436 546500 14464
rect 414072 14424 414078 14436
rect 546494 14424 546500 14436
rect 546552 14424 546558 14476
rect 280154 13676 280160 13728
rect 280212 13716 280218 13728
rect 392486 13716 392492 13728
rect 280212 13688 392492 13716
rect 280212 13676 280218 13688
rect 392486 13676 392492 13688
rect 392544 13676 392550 13728
rect 281534 13608 281540 13660
rect 281592 13648 281598 13660
rect 396166 13648 396172 13660
rect 281592 13620 396172 13648
rect 281592 13608 281598 13620
rect 396166 13608 396172 13620
rect 396224 13608 396230 13660
rect 281626 13540 281632 13592
rect 281684 13580 281690 13592
rect 400122 13580 400128 13592
rect 281684 13552 400128 13580
rect 281684 13540 281690 13552
rect 400122 13540 400128 13552
rect 400180 13540 400186 13592
rect 217318 13472 217324 13524
rect 217376 13512 217382 13524
rect 242894 13512 242900 13524
rect 217376 13484 242900 13512
rect 217376 13472 217382 13484
rect 242894 13472 242900 13484
rect 242952 13472 242958 13524
rect 282914 13472 282920 13524
rect 282972 13512 282978 13524
rect 403618 13512 403624 13524
rect 282972 13484 403624 13512
rect 282972 13472 282978 13484
rect 403618 13472 403624 13484
rect 403676 13472 403682 13524
rect 404354 13472 404360 13524
rect 404412 13512 404418 13524
rect 503714 13512 503720 13524
rect 404412 13484 503720 13512
rect 404412 13472 404418 13484
rect 503714 13472 503720 13484
rect 503772 13472 503778 13524
rect 215294 13404 215300 13456
rect 215352 13444 215358 13456
rect 241514 13444 241520 13456
rect 215352 13416 241520 13444
rect 215352 13404 215358 13416
rect 241514 13404 241520 13416
rect 241572 13404 241578 13456
rect 284386 13404 284392 13456
rect 284444 13444 284450 13456
rect 407114 13444 407120 13456
rect 284444 13416 407120 13444
rect 284444 13404 284450 13416
rect 407114 13404 407120 13416
rect 407172 13404 407178 13456
rect 132586 13336 132592 13388
rect 132644 13376 132650 13388
rect 175458 13376 175464 13388
rect 132644 13348 175464 13376
rect 132644 13336 132650 13348
rect 175458 13336 175464 13348
rect 175516 13336 175522 13388
rect 201586 13336 201592 13388
rect 201644 13376 201650 13388
rect 238754 13376 238760 13388
rect 201644 13348 238760 13376
rect 201644 13336 201650 13348
rect 238754 13336 238760 13348
rect 238812 13336 238818 13388
rect 284294 13336 284300 13388
rect 284352 13376 284358 13388
rect 410794 13376 410800 13388
rect 284352 13348 410800 13376
rect 284352 13336 284358 13348
rect 410794 13336 410800 13348
rect 410852 13336 410858 13388
rect 411254 13336 411260 13388
rect 411312 13376 411318 13388
rect 536098 13376 536104 13388
rect 411312 13348 536104 13376
rect 411312 13336 411318 13348
rect 536098 13336 536104 13348
rect 536156 13336 536162 13388
rect 166074 13268 166080 13320
rect 166132 13308 166138 13320
rect 230474 13308 230480 13320
rect 166132 13280 230480 13308
rect 166132 13268 166138 13280
rect 230474 13268 230480 13280
rect 230532 13268 230538 13320
rect 285766 13268 285772 13320
rect 285824 13308 285830 13320
rect 417418 13308 417424 13320
rect 285824 13280 417424 13308
rect 285824 13268 285830 13280
rect 417418 13268 417424 13280
rect 417476 13268 417482 13320
rect 154666 13200 154672 13252
rect 154724 13240 154730 13252
rect 274818 13240 274824 13252
rect 154724 13212 274824 13240
rect 154724 13200 154730 13212
rect 274818 13200 274824 13212
rect 274876 13200 274882 13252
rect 287146 13200 287152 13252
rect 287204 13240 287210 13252
rect 421006 13240 421012 13252
rect 287204 13212 421012 13240
rect 287204 13200 287210 13212
rect 421006 13200 421012 13212
rect 421064 13200 421070 13252
rect 63494 13132 63500 13184
rect 63552 13172 63558 13184
rect 111610 13172 111616 13184
rect 63552 13144 111616 13172
rect 63552 13132 63558 13144
rect 111610 13132 111616 13144
rect 111668 13132 111674 13184
rect 163682 13132 163688 13184
rect 163740 13172 163746 13184
rect 286318 13172 286324 13184
rect 163740 13144 286324 13172
rect 163740 13132 163746 13144
rect 286318 13132 286324 13144
rect 286376 13132 286382 13184
rect 287054 13132 287060 13184
rect 287112 13172 287118 13184
rect 424962 13172 424968 13184
rect 287112 13144 424968 13172
rect 287112 13132 287118 13144
rect 424962 13132 424968 13144
rect 425020 13132 425026 13184
rect 30098 13064 30104 13116
rect 30156 13104 30162 13116
rect 45554 13104 45560 13116
rect 30156 13076 45560 13104
rect 30156 13064 30162 13076
rect 45554 13064 45560 13076
rect 45612 13064 45618 13116
rect 53282 13064 53288 13116
rect 53340 13104 53346 13116
rect 100754 13104 100760 13116
rect 53340 13076 100760 13104
rect 53340 13064 53346 13076
rect 100754 13064 100760 13076
rect 100812 13064 100818 13116
rect 138842 13064 138848 13116
rect 138900 13104 138906 13116
rect 282178 13104 282184 13116
rect 138900 13076 282184 13104
rect 138900 13064 138906 13076
rect 282178 13064 282184 13076
rect 282236 13064 282242 13116
rect 285674 13064 285680 13116
rect 285732 13104 285738 13116
rect 414290 13104 414296 13116
rect 285732 13076 414296 13104
rect 285732 13064 285738 13076
rect 414290 13064 414296 13076
rect 414348 13064 414354 13116
rect 414658 13064 414664 13116
rect 414716 13104 414722 13116
rect 576946 13104 576952 13116
rect 414716 13076 576952 13104
rect 414716 13064 414722 13076
rect 576946 13064 576952 13076
rect 577004 13064 577010 13116
rect 249886 12316 249892 12368
rect 249944 12356 249950 12368
rect 254210 12356 254216 12368
rect 249944 12328 254216 12356
rect 249944 12316 249950 12328
rect 254210 12316 254216 12328
rect 254268 12316 254274 12368
rect 197906 12248 197912 12300
rect 197964 12288 197970 12300
rect 237374 12288 237380 12300
rect 197964 12260 237380 12288
rect 197964 12248 197970 12260
rect 237374 12248 237380 12260
rect 237432 12248 237438 12300
rect 266446 12248 266452 12300
rect 266504 12288 266510 12300
rect 324406 12288 324412 12300
rect 266504 12260 324412 12288
rect 266504 12248 266510 12260
rect 324406 12248 324412 12260
rect 324464 12248 324470 12300
rect 190638 12180 190644 12232
rect 190696 12220 190702 12232
rect 235994 12220 236000 12232
rect 190696 12192 236000 12220
rect 190696 12180 190702 12192
rect 235994 12180 236000 12192
rect 236052 12180 236058 12232
rect 266354 12180 266360 12232
rect 266412 12220 266418 12232
rect 328730 12220 328736 12232
rect 266412 12192 328736 12220
rect 266412 12180 266418 12192
rect 328730 12180 328736 12192
rect 328788 12180 328794 12232
rect 186866 12112 186872 12164
rect 186924 12152 186930 12164
rect 234706 12152 234712 12164
rect 186924 12124 234712 12152
rect 186924 12112 186930 12124
rect 234706 12112 234712 12124
rect 234764 12112 234770 12164
rect 267734 12112 267740 12164
rect 267792 12152 267798 12164
rect 336274 12152 336280 12164
rect 267792 12124 336280 12152
rect 267792 12112 267798 12124
rect 336274 12112 336280 12124
rect 336332 12112 336338 12164
rect 183738 12044 183744 12096
rect 183796 12084 183802 12096
rect 234798 12084 234804 12096
rect 183796 12056 234804 12084
rect 183796 12044 183802 12056
rect 234798 12044 234804 12056
rect 234856 12044 234862 12096
rect 269206 12044 269212 12096
rect 269264 12084 269270 12096
rect 339494 12084 339500 12096
rect 269264 12056 339500 12084
rect 269264 12044 269270 12056
rect 339494 12044 339500 12056
rect 339552 12044 339558 12096
rect 180242 11976 180248 12028
rect 180300 12016 180306 12028
rect 233326 12016 233332 12028
rect 180300 11988 233332 12016
rect 180300 11976 180306 11988
rect 233326 11976 233332 11988
rect 233384 11976 233390 12028
rect 269114 11976 269120 12028
rect 269172 12016 269178 12028
rect 342898 12016 342904 12028
rect 269172 11988 342904 12016
rect 269172 11976 269178 11988
rect 342898 11976 342904 11988
rect 342956 11976 342962 12028
rect 393958 11976 393964 12028
rect 394016 12016 394022 12028
rect 415486 12016 415492 12028
rect 394016 11988 415492 12016
rect 394016 11976 394022 11988
rect 415486 11976 415492 11988
rect 415544 11976 415550 12028
rect 176838 11908 176844 11960
rect 176896 11948 176902 11960
rect 233234 11948 233240 11960
rect 176896 11920 233240 11948
rect 176896 11908 176902 11920
rect 233234 11908 233240 11920
rect 233292 11908 233298 11960
rect 270586 11908 270592 11960
rect 270644 11948 270650 11960
rect 346946 11948 346952 11960
rect 270644 11920 346952 11948
rect 270644 11908 270650 11920
rect 346946 11908 346952 11920
rect 347004 11908 347010 11960
rect 383654 11908 383660 11960
rect 383712 11948 383718 11960
rect 407206 11948 407212 11960
rect 383712 11920 407212 11948
rect 383712 11908 383718 11920
rect 407206 11908 407212 11920
rect 407264 11908 407270 11960
rect 172698 11840 172704 11892
rect 172756 11880 172762 11892
rect 231946 11880 231952 11892
rect 172756 11852 231952 11880
rect 172756 11840 172762 11852
rect 231946 11840 231952 11852
rect 232004 11840 232010 11892
rect 249794 11840 249800 11892
rect 249852 11880 249858 11892
rect 251450 11880 251456 11892
rect 249852 11852 251456 11880
rect 249852 11840 249858 11852
rect 251450 11840 251456 11852
rect 251508 11840 251514 11892
rect 271874 11840 271880 11892
rect 271932 11880 271938 11892
rect 353570 11880 353576 11892
rect 271932 11852 353576 11880
rect 271932 11840 271938 11852
rect 353570 11840 353576 11852
rect 353628 11840 353634 11892
rect 405826 11840 405832 11892
rect 405884 11880 405890 11892
rect 511258 11880 511264 11892
rect 405884 11852 511264 11880
rect 405884 11840 405890 11852
rect 511258 11840 511264 11852
rect 511316 11840 511322 11892
rect 37826 11772 37832 11824
rect 37884 11812 37890 11824
rect 71038 11812 71044 11824
rect 37884 11784 71044 11812
rect 37884 11772 37890 11784
rect 71038 11772 71044 11784
rect 71096 11772 71102 11824
rect 85666 11772 85672 11824
rect 85724 11812 85730 11824
rect 107654 11812 107660 11824
rect 85724 11784 107660 11812
rect 85724 11772 85730 11784
rect 107654 11772 107660 11784
rect 107712 11772 107718 11824
rect 168374 11772 168380 11824
rect 168432 11812 168438 11824
rect 231854 11812 231860 11824
rect 168432 11784 231860 11812
rect 168432 11772 168438 11784
rect 231854 11772 231860 11784
rect 231912 11772 231918 11824
rect 236546 11772 236552 11824
rect 236604 11812 236610 11824
rect 245746 11812 245752 11824
rect 236604 11784 245752 11812
rect 236604 11772 236610 11784
rect 245746 11772 245752 11784
rect 245804 11772 245810 11824
rect 270678 11772 270684 11824
rect 270736 11812 270742 11824
rect 349246 11812 349252 11824
rect 270736 11784 349252 11812
rect 270736 11772 270742 11784
rect 349246 11772 349252 11784
rect 349304 11772 349310 11824
rect 349798 11772 349804 11824
rect 349856 11812 349862 11824
rect 531314 11812 531320 11824
rect 349856 11784 531320 11812
rect 349856 11772 349862 11784
rect 531314 11772 531320 11784
rect 531372 11772 531378 11824
rect 60826 11704 60832 11756
rect 60884 11744 60890 11756
rect 100754 11744 100760 11756
rect 60884 11716 100760 11744
rect 60884 11704 60890 11716
rect 100754 11704 100760 11716
rect 100812 11704 100818 11756
rect 105538 11704 105544 11756
rect 105596 11744 105602 11756
rect 119890 11744 119896 11756
rect 105596 11716 119896 11744
rect 105596 11704 105602 11716
rect 119890 11704 119896 11716
rect 119948 11704 119954 11756
rect 130562 11704 130568 11756
rect 130620 11744 130626 11756
rect 222286 11744 222292 11756
rect 130620 11716 222292 11744
rect 130620 11704 130626 11716
rect 222286 11704 222292 11716
rect 222344 11704 222350 11756
rect 233418 11704 233424 11756
rect 233476 11744 233482 11756
rect 244918 11744 244924 11756
rect 233476 11716 244924 11744
rect 233476 11704 233482 11716
rect 244918 11704 244924 11716
rect 244976 11704 244982 11756
rect 273346 11704 273352 11756
rect 273404 11744 273410 11756
rect 357526 11744 357532 11756
rect 273404 11716 357532 11744
rect 273404 11704 273410 11716
rect 357526 11704 357532 11716
rect 357584 11704 357590 11756
rect 360838 11704 360844 11756
rect 360896 11744 360902 11756
rect 562042 11744 562048 11756
rect 360896 11716 562048 11744
rect 360896 11704 360902 11716
rect 562042 11704 562048 11716
rect 562100 11704 562106 11756
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 423674 11568 423680 11620
rect 423732 11608 423738 11620
rect 423732 11580 423812 11608
rect 423732 11568 423738 11580
rect 423784 11416 423812 11580
rect 240226 11364 240232 11416
rect 240284 11404 240290 11416
rect 247034 11404 247040 11416
rect 240284 11376 247040 11404
rect 240284 11364 240290 11376
rect 247034 11364 247040 11376
rect 247092 11364 247098 11416
rect 423766 11364 423772 11416
rect 423824 11364 423830 11416
rect 187694 10616 187700 10668
rect 187752 10656 187758 10668
rect 423858 10656 423864 10668
rect 187752 10628 423864 10656
rect 187752 10616 187758 10628
rect 423858 10616 423864 10628
rect 423916 10616 423922 10668
rect 425698 10616 425704 10668
rect 425756 10656 425762 10668
rect 532050 10656 532056 10668
rect 425756 10628 532056 10656
rect 425756 10616 425762 10628
rect 532050 10616 532056 10628
rect 532108 10616 532114 10668
rect 190546 10548 190552 10600
rect 190604 10588 190610 10600
rect 433978 10588 433984 10600
rect 190604 10560 433984 10588
rect 190604 10548 190610 10560
rect 433978 10548 433984 10560
rect 434036 10548 434042 10600
rect 436738 10548 436744 10600
rect 436796 10588 436802 10600
rect 550266 10588 550272 10600
rect 436796 10560 550272 10588
rect 436796 10548 436802 10560
rect 550266 10548 550272 10560
rect 550324 10548 550330 10600
rect 190454 10480 190460 10532
rect 190512 10520 190518 10532
rect 437474 10520 437480 10532
rect 190512 10492 437480 10520
rect 190512 10480 190518 10492
rect 437474 10480 437480 10492
rect 437532 10480 437538 10532
rect 191926 10412 191932 10464
rect 191984 10452 191990 10464
rect 440326 10452 440332 10464
rect 191984 10424 440332 10452
rect 191984 10412 191990 10424
rect 440326 10412 440332 10424
rect 440384 10412 440390 10464
rect 41874 10344 41880 10396
rect 41932 10384 41938 10396
rect 72418 10384 72424 10396
rect 41932 10356 72424 10384
rect 41932 10344 41938 10356
rect 72418 10344 72424 10356
rect 72476 10344 72482 10396
rect 89714 10344 89720 10396
rect 89772 10384 89778 10396
rect 112346 10384 112352 10396
rect 89772 10356 112352 10384
rect 89772 10344 89778 10356
rect 112346 10344 112352 10356
rect 112404 10344 112410 10396
rect 191834 10344 191840 10396
rect 191892 10384 191898 10396
rect 445018 10384 445024 10396
rect 191892 10356 445024 10384
rect 191892 10344 191898 10356
rect 445018 10344 445024 10356
rect 445076 10344 445082 10396
rect 17034 10276 17040 10328
rect 17092 10316 17098 10328
rect 42794 10316 42800 10328
rect 17092 10288 42800 10316
rect 17092 10276 17098 10288
rect 42794 10276 42800 10288
rect 42852 10276 42858 10328
rect 60734 10276 60740 10328
rect 60792 10316 60798 10328
rect 97442 10316 97448 10328
rect 60792 10288 97448 10316
rect 60792 10276 60798 10288
rect 97442 10276 97448 10288
rect 97500 10276 97506 10328
rect 132494 10276 132500 10328
rect 132552 10316 132558 10328
rect 171962 10316 171968 10328
rect 132552 10288 171968 10316
rect 132552 10276 132558 10288
rect 171962 10276 171968 10288
rect 172020 10276 172026 10328
rect 177298 10276 177304 10328
rect 177356 10316 177362 10328
rect 186130 10316 186136 10328
rect 177356 10288 186136 10316
rect 177356 10276 177362 10288
rect 186130 10276 186136 10288
rect 186188 10276 186194 10328
rect 194594 10276 194600 10328
rect 194652 10316 194658 10328
rect 455690 10316 455696 10328
rect 194652 10288 455696 10316
rect 194652 10276 194658 10288
rect 455690 10276 455696 10288
rect 455748 10276 455754 10328
rect 172514 9528 172520 9580
rect 172572 9568 172578 9580
rect 356330 9568 356336 9580
rect 172572 9540 356336 9568
rect 172572 9528 172578 9540
rect 356330 9528 356336 9540
rect 356388 9528 356394 9580
rect 173986 9460 173992 9512
rect 174044 9500 174050 9512
rect 359918 9500 359924 9512
rect 174044 9472 359924 9500
rect 174044 9460 174050 9472
rect 359918 9460 359924 9472
rect 359976 9460 359982 9512
rect 173894 9392 173900 9444
rect 173952 9432 173958 9444
rect 363506 9432 363512 9444
rect 173952 9404 363512 9432
rect 173952 9392 173958 9404
rect 363506 9392 363512 9404
rect 363564 9392 363570 9444
rect 175274 9324 175280 9376
rect 175332 9364 175338 9376
rect 367002 9364 367008 9376
rect 175332 9336 367008 9364
rect 175332 9324 175338 9336
rect 367002 9324 367008 9336
rect 367060 9324 367066 9376
rect 175366 9256 175372 9308
rect 175424 9296 175430 9308
rect 370590 9296 370596 9308
rect 175424 9268 370596 9296
rect 175424 9256 175430 9268
rect 370590 9256 370596 9268
rect 370648 9256 370654 9308
rect 382274 9256 382280 9308
rect 382332 9296 382338 9308
rect 404814 9296 404820 9308
rect 382332 9268 404820 9296
rect 382332 9256 382338 9268
rect 404814 9256 404820 9268
rect 404872 9256 404878 9308
rect 176654 9188 176660 9240
rect 176712 9228 176718 9240
rect 374086 9228 374092 9240
rect 176712 9200 374092 9228
rect 176712 9188 176718 9200
rect 374086 9188 374092 9200
rect 374144 9188 374150 9240
rect 380986 9188 380992 9240
rect 381044 9228 381050 9240
rect 397730 9228 397736 9240
rect 381044 9200 397736 9228
rect 381044 9188 381050 9200
rect 397730 9188 397736 9200
rect 397788 9188 397794 9240
rect 400214 9188 400220 9240
rect 400272 9228 400278 9240
rect 482830 9228 482836 9240
rect 400272 9200 482836 9228
rect 400272 9188 400278 9200
rect 482830 9188 482836 9200
rect 482888 9188 482894 9240
rect 178034 9120 178040 9172
rect 178092 9160 178098 9172
rect 377674 9160 377680 9172
rect 178092 9132 377680 9160
rect 178092 9120 178098 9132
rect 377674 9120 377680 9132
rect 377732 9120 377738 9172
rect 400306 9120 400312 9172
rect 400364 9160 400370 9172
rect 486418 9160 486424 9172
rect 400364 9132 486424 9160
rect 400364 9120 400370 9132
rect 486418 9120 486424 9132
rect 486476 9120 486482 9172
rect 85758 9052 85764 9104
rect 85816 9092 85822 9104
rect 95142 9092 95148 9104
rect 85816 9064 95148 9092
rect 85816 9052 85822 9064
rect 95142 9052 95148 9064
rect 95200 9052 95206 9104
rect 178126 9052 178132 9104
rect 178184 9092 178190 9104
rect 381170 9092 381176 9104
rect 178184 9064 381176 9092
rect 178184 9052 178190 9064
rect 381170 9052 381176 9064
rect 381228 9052 381234 9104
rect 401594 9052 401600 9104
rect 401652 9092 401658 9104
rect 489914 9092 489920 9104
rect 401652 9064 489920 9092
rect 401652 9052 401658 9064
rect 489914 9052 489920 9064
rect 489972 9052 489978 9104
rect 53926 8984 53932 9036
rect 53984 9024 53990 9036
rect 69106 9024 69112 9036
rect 53984 8996 69112 9024
rect 53984 8984 53990 8996
rect 69106 8984 69112 8996
rect 69164 8984 69170 9036
rect 70302 8984 70308 9036
rect 70360 9024 70366 9036
rect 80146 9024 80152 9036
rect 70360 8996 80152 9024
rect 70360 8984 70366 8996
rect 80146 8984 80152 8996
rect 80204 8984 80210 9036
rect 87046 8984 87052 9036
rect 87104 9024 87110 9036
rect 102226 9024 102232 9036
rect 87104 8996 102232 9024
rect 87104 8984 87110 8996
rect 102226 8984 102232 8996
rect 102284 8984 102290 9036
rect 146938 8984 146944 9036
rect 146996 9024 147002 9036
rect 168466 9024 168472 9036
rect 146996 8996 168472 9024
rect 146996 8984 147002 8996
rect 168466 8984 168472 8996
rect 168524 8984 168530 9036
rect 179414 8984 179420 9036
rect 179472 9024 179478 9036
rect 384758 9024 384764 9036
rect 179472 8996 384764 9024
rect 179472 8984 179478 8996
rect 384758 8984 384764 8996
rect 384816 8984 384822 9036
rect 403066 8984 403072 9036
rect 403124 9024 403130 9036
rect 493502 9024 493508 9036
rect 403124 8996 493508 9024
rect 403124 8984 403130 8996
rect 493502 8984 493508 8996
rect 493560 8984 493566 9036
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 40126 8956 40132 8968
rect 4028 8928 40132 8956
rect 4028 8916 4034 8928
rect 40126 8916 40132 8928
rect 40184 8916 40190 8968
rect 63218 8916 63224 8968
rect 63276 8956 63282 8968
rect 78674 8956 78680 8968
rect 63276 8928 78680 8956
rect 63276 8916 63282 8928
rect 78674 8916 78680 8928
rect 78732 8916 78738 8968
rect 93118 8916 93124 8968
rect 93176 8956 93182 8968
rect 116394 8956 116400 8968
rect 93176 8928 116400 8956
rect 93176 8916 93182 8928
rect 116394 8916 116400 8928
rect 116452 8916 116458 8968
rect 128354 8916 128360 8968
rect 128412 8956 128418 8968
rect 154206 8956 154212 8968
rect 128412 8928 154212 8956
rect 128412 8916 128418 8928
rect 154206 8916 154212 8928
rect 154264 8916 154270 8968
rect 179506 8916 179512 8968
rect 179564 8956 179570 8968
rect 388254 8956 388260 8968
rect 179564 8928 388260 8956
rect 179564 8916 179570 8928
rect 388254 8916 388260 8928
rect 388312 8916 388318 8968
rect 392578 8916 392584 8968
rect 392636 8956 392642 8968
rect 401318 8956 401324 8968
rect 392636 8928 401324 8956
rect 392636 8916 392642 8928
rect 401318 8916 401324 8928
rect 401376 8916 401382 8968
rect 402974 8916 402980 8968
rect 403032 8956 403038 8968
rect 497090 8956 497096 8968
rect 403032 8928 497096 8956
rect 403032 8916 403038 8928
rect 497090 8916 497096 8928
rect 497148 8916 497154 8968
rect 80882 8712 80888 8764
rect 80940 8752 80946 8764
rect 82906 8752 82912 8764
rect 80940 8724 82912 8752
rect 80940 8712 80946 8724
rect 82906 8712 82912 8724
rect 82964 8712 82970 8764
rect 284294 8168 284300 8220
rect 284352 8208 284358 8220
rect 324958 8208 324964 8220
rect 284352 8180 324964 8208
rect 284352 8168 284358 8180
rect 324958 8168 324964 8180
rect 325016 8168 325022 8220
rect 263594 8100 263600 8152
rect 263652 8140 263658 8152
rect 318518 8140 318524 8152
rect 263652 8112 318524 8140
rect 263652 8100 263658 8112
rect 318518 8100 318524 8112
rect 318576 8100 318582 8152
rect 131758 8032 131764 8084
rect 131816 8072 131822 8084
rect 322198 8072 322204 8084
rect 131816 8044 322204 8072
rect 131816 8032 131822 8044
rect 322198 8032 322204 8044
rect 322256 8032 322262 8084
rect 313366 7964 313372 8016
rect 313424 8004 313430 8016
rect 541986 8004 541992 8016
rect 313424 7976 541992 8004
rect 313424 7964 313430 7976
rect 541986 7964 541992 7976
rect 542044 7964 542050 8016
rect 316034 7896 316040 7948
rect 316092 7936 316098 7948
rect 552658 7936 552664 7948
rect 316092 7908 552664 7936
rect 316092 7896 316098 7908
rect 552658 7896 552664 7908
rect 552716 7896 552722 7948
rect 316126 7828 316132 7880
rect 316184 7868 316190 7880
rect 556154 7868 556160 7880
rect 316184 7840 556160 7868
rect 316184 7828 316190 7840
rect 556154 7828 556160 7840
rect 556212 7828 556218 7880
rect 208578 7760 208584 7812
rect 208636 7800 208642 7812
rect 240134 7800 240140 7812
rect 208636 7772 240140 7800
rect 208636 7760 208642 7772
rect 240134 7760 240140 7772
rect 240192 7760 240198 7812
rect 259546 7760 259552 7812
rect 259604 7800 259610 7812
rect 297266 7800 297272 7812
rect 259604 7772 297272 7800
rect 259604 7760 259610 7772
rect 297266 7760 297272 7772
rect 297324 7760 297330 7812
rect 317414 7760 317420 7812
rect 317472 7800 317478 7812
rect 559742 7800 559748 7812
rect 317472 7772 559748 7800
rect 317472 7760 317478 7772
rect 559742 7760 559748 7772
rect 559800 7760 559806 7812
rect 85574 7692 85580 7744
rect 85632 7732 85638 7744
rect 98638 7732 98644 7744
rect 85632 7704 98644 7732
rect 85632 7692 85638 7704
rect 98638 7692 98644 7704
rect 98696 7692 98702 7744
rect 160094 7692 160100 7744
rect 160152 7732 160158 7744
rect 299658 7732 299664 7744
rect 160152 7704 299664 7732
rect 160152 7692 160158 7704
rect 299658 7692 299664 7704
rect 299716 7692 299722 7744
rect 317506 7692 317512 7744
rect 317564 7732 317570 7744
rect 563238 7732 563244 7744
rect 317564 7704 563244 7732
rect 317564 7692 317570 7704
rect 563238 7692 563244 7704
rect 563296 7692 563302 7744
rect 53834 7624 53840 7676
rect 53892 7664 53898 7676
rect 65518 7664 65524 7676
rect 53892 7636 65524 7664
rect 53892 7624 53898 7636
rect 65518 7624 65524 7636
rect 65576 7624 65582 7676
rect 69658 7624 69664 7676
rect 69716 7664 69722 7676
rect 90358 7664 90364 7676
rect 69716 7636 90364 7664
rect 69716 7624 69722 7636
rect 90358 7624 90364 7636
rect 90416 7624 90422 7676
rect 161658 7624 161664 7676
rect 161716 7664 161722 7676
rect 303154 7664 303160 7676
rect 161716 7636 303160 7664
rect 161716 7624 161722 7636
rect 303154 7624 303160 7636
rect 303212 7624 303218 7676
rect 320266 7624 320272 7676
rect 320324 7664 320330 7676
rect 570322 7664 570328 7676
rect 320324 7636 570328 7664
rect 320324 7624 320330 7636
rect 570322 7624 570328 7636
rect 570380 7624 570386 7676
rect 26510 7556 26516 7608
rect 26568 7596 26574 7608
rect 44174 7596 44180 7608
rect 26568 7568 44180 7596
rect 26568 7556 26574 7568
rect 44174 7556 44180 7568
rect 44232 7556 44238 7608
rect 59630 7556 59636 7608
rect 59688 7596 59694 7608
rect 75178 7596 75184 7608
rect 59688 7568 75184 7596
rect 59688 7556 59694 7568
rect 75178 7556 75184 7568
rect 75236 7556 75242 7608
rect 88334 7556 88340 7608
rect 88392 7596 88398 7608
rect 109310 7596 109316 7608
rect 88392 7568 109316 7596
rect 88392 7556 88398 7568
rect 109310 7556 109316 7568
rect 109368 7556 109374 7608
rect 141418 7556 141424 7608
rect 141476 7596 141482 7608
rect 161290 7596 161296 7608
rect 141476 7568 161296 7596
rect 141476 7556 141482 7568
rect 161290 7556 161296 7568
rect 161348 7556 161354 7608
rect 161566 7556 161572 7608
rect 161624 7596 161630 7608
rect 306742 7596 306748 7608
rect 161624 7568 306748 7596
rect 161624 7556 161630 7568
rect 306742 7556 306748 7568
rect 306800 7556 306806 7608
rect 320174 7556 320180 7608
rect 320232 7596 320238 7608
rect 573910 7596 573916 7608
rect 320232 7568 573916 7596
rect 320232 7556 320238 7568
rect 573910 7556 573916 7568
rect 573968 7556 573974 7608
rect 218054 7488 218060 7540
rect 218112 7528 218118 7540
rect 219250 7528 219256 7540
rect 218112 7500 219256 7528
rect 218112 7488 218118 7500
rect 219250 7488 219256 7500
rect 219308 7488 219314 7540
rect 77386 7216 77392 7268
rect 77444 7256 77450 7268
rect 81434 7256 81440 7268
rect 77444 7228 81440 7256
rect 77444 7216 77450 7228
rect 81434 7216 81440 7228
rect 81492 7216 81498 7268
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 37918 6848 37924 6860
rect 3476 6820 37924 6848
rect 3476 6808 3482 6820
rect 37918 6808 37924 6820
rect 37976 6808 37982 6860
rect 252646 6808 252652 6860
rect 252704 6848 252710 6860
rect 265342 6848 265348 6860
rect 252704 6820 265348 6848
rect 252704 6808 252710 6820
rect 265342 6808 265348 6820
rect 265400 6808 265406 6860
rect 428550 6808 428556 6860
rect 428608 6848 428614 6860
rect 580166 6848 580172 6860
rect 428608 6820 580172 6848
rect 428608 6808 428614 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 264974 6672 264980 6724
rect 265032 6712 265038 6724
rect 322106 6712 322112 6724
rect 265032 6684 322112 6712
rect 265032 6672 265038 6684
rect 322106 6672 322112 6684
rect 322164 6672 322170 6724
rect 251358 6604 251364 6656
rect 251416 6644 251422 6656
rect 261754 6644 261760 6656
rect 251416 6616 261760 6644
rect 251416 6604 251422 6616
rect 261754 6604 261760 6616
rect 261812 6604 261818 6656
rect 299474 6604 299480 6656
rect 299532 6644 299538 6656
rect 481726 6644 481732 6656
rect 299532 6616 481732 6644
rect 299532 6604 299538 6616
rect 481726 6604 481732 6616
rect 481784 6604 481790 6656
rect 252554 6536 252560 6588
rect 252612 6576 252618 6588
rect 268838 6576 268844 6588
rect 252612 6548 268844 6576
rect 252612 6536 252618 6548
rect 268838 6536 268844 6548
rect 268896 6536 268902 6588
rect 300854 6536 300860 6588
rect 300912 6576 300918 6588
rect 485222 6576 485228 6588
rect 300912 6548 485228 6576
rect 300912 6536 300918 6548
rect 485222 6536 485228 6548
rect 485280 6536 485286 6588
rect 143534 6468 143540 6520
rect 143592 6508 143598 6520
rect 225138 6508 225144 6520
rect 143592 6480 225144 6508
rect 143592 6468 143598 6480
rect 225138 6468 225144 6480
rect 225196 6468 225202 6520
rect 253934 6468 253940 6520
rect 253992 6508 253998 6520
rect 272426 6508 272432 6520
rect 253992 6480 272432 6508
rect 253992 6468 253998 6480
rect 272426 6468 272432 6480
rect 272484 6468 272490 6520
rect 302234 6468 302240 6520
rect 302292 6508 302298 6520
rect 488810 6508 488816 6520
rect 302292 6480 488816 6508
rect 302292 6468 302298 6480
rect 488810 6468 488816 6480
rect 488868 6468 488874 6520
rect 144914 6400 144920 6452
rect 144972 6440 144978 6452
rect 228726 6440 228732 6452
rect 144972 6412 228732 6440
rect 144972 6400 144978 6412
rect 228726 6400 228732 6412
rect 228784 6400 228790 6452
rect 229830 6400 229836 6452
rect 229888 6440 229894 6452
rect 244458 6440 244464 6452
rect 229888 6412 244464 6440
rect 229888 6400 229894 6412
rect 244458 6400 244464 6412
rect 244516 6400 244522 6452
rect 255406 6400 255412 6452
rect 255464 6440 255470 6452
rect 276014 6440 276020 6452
rect 255464 6412 276020 6440
rect 255464 6400 255470 6412
rect 276014 6400 276020 6412
rect 276072 6400 276078 6452
rect 302326 6400 302332 6452
rect 302384 6440 302390 6452
rect 492306 6440 492312 6452
rect 302384 6412 492312 6440
rect 302384 6400 302390 6412
rect 492306 6400 492312 6412
rect 492364 6400 492370 6452
rect 145006 6332 145012 6384
rect 145064 6372 145070 6384
rect 232222 6372 232228 6384
rect 145064 6344 232228 6372
rect 145064 6332 145070 6344
rect 232222 6332 232228 6344
rect 232280 6332 232286 6384
rect 255314 6332 255320 6384
rect 255372 6372 255378 6384
rect 279510 6372 279516 6384
rect 255372 6344 279516 6372
rect 255372 6332 255378 6344
rect 279510 6332 279516 6344
rect 279568 6332 279574 6384
rect 303798 6332 303804 6384
rect 303856 6372 303862 6384
rect 495894 6372 495900 6384
rect 303856 6344 495900 6372
rect 303856 6332 303862 6344
rect 495894 6332 495900 6344
rect 495952 6332 495958 6384
rect 146294 6264 146300 6316
rect 146352 6304 146358 6316
rect 235810 6304 235816 6316
rect 146352 6276 235816 6304
rect 146352 6264 146358 6276
rect 235810 6264 235816 6276
rect 235868 6264 235874 6316
rect 256694 6264 256700 6316
rect 256752 6304 256758 6316
rect 283098 6304 283104 6316
rect 256752 6276 283104 6304
rect 256752 6264 256758 6276
rect 283098 6264 283104 6276
rect 283156 6264 283162 6316
rect 303706 6264 303712 6316
rect 303764 6304 303770 6316
rect 499390 6304 499396 6316
rect 303764 6276 499396 6304
rect 303764 6264 303770 6276
rect 499390 6264 499396 6276
rect 499448 6264 499454 6316
rect 58618 6196 58624 6248
rect 58676 6236 58682 6248
rect 72602 6236 72608 6248
rect 58676 6208 72608 6236
rect 58676 6196 58682 6208
rect 72602 6196 72608 6208
rect 72660 6196 72666 6248
rect 73798 6196 73804 6248
rect 73856 6236 73862 6248
rect 80054 6236 80060 6248
rect 73856 6208 80060 6236
rect 73856 6196 73862 6208
rect 80054 6196 80060 6208
rect 80112 6196 80118 6248
rect 147674 6196 147680 6248
rect 147732 6236 147738 6248
rect 239306 6236 239312 6248
rect 147732 6208 239312 6236
rect 147732 6196 147738 6208
rect 239306 6196 239312 6208
rect 239364 6196 239370 6248
rect 256786 6196 256792 6248
rect 256844 6236 256850 6248
rect 286594 6236 286600 6248
rect 256844 6208 286600 6236
rect 256844 6196 256850 6208
rect 286594 6196 286600 6208
rect 286652 6196 286658 6248
rect 304994 6196 305000 6248
rect 305052 6236 305058 6248
rect 502978 6236 502984 6248
rect 305052 6208 502984 6236
rect 305052 6196 305058 6208
rect 502978 6196 502984 6208
rect 503036 6196 503042 6248
rect 52546 6128 52552 6180
rect 52604 6168 52610 6180
rect 58434 6168 58440 6180
rect 52604 6140 58440 6168
rect 52604 6128 52610 6140
rect 58434 6128 58440 6140
rect 58492 6128 58498 6180
rect 64874 6128 64880 6180
rect 64932 6168 64938 6180
rect 118786 6168 118792 6180
rect 64932 6140 118792 6168
rect 64932 6128 64938 6140
rect 118786 6128 118792 6140
rect 118844 6128 118850 6180
rect 150434 6128 150440 6180
rect 150492 6168 150498 6180
rect 253474 6168 253480 6180
rect 150492 6140 253480 6168
rect 150492 6128 150498 6140
rect 253474 6128 253480 6140
rect 253532 6128 253538 6180
rect 258166 6128 258172 6180
rect 258224 6168 258230 6180
rect 293678 6168 293684 6180
rect 258224 6140 293684 6168
rect 258224 6128 258230 6140
rect 293678 6128 293684 6140
rect 293736 6128 293742 6180
rect 305086 6128 305092 6180
rect 305144 6168 305150 6180
rect 506474 6168 506480 6180
rect 305144 6140 506480 6168
rect 305144 6128 305150 6140
rect 506474 6128 506480 6140
rect 506532 6128 506538 6180
rect 244090 5584 244096 5636
rect 244148 5624 244154 5636
rect 248506 5624 248512 5636
rect 244148 5596 248512 5624
rect 244148 5584 244154 5596
rect 248506 5584 248512 5596
rect 248564 5584 248570 5636
rect 44266 5516 44272 5568
rect 44324 5556 44330 5568
rect 46198 5556 46204 5568
rect 44324 5528 46204 5556
rect 44324 5516 44330 5528
rect 46198 5516 46204 5528
rect 46256 5516 46262 5568
rect 84194 5516 84200 5568
rect 84252 5556 84258 5568
rect 91554 5556 91560 5568
rect 84252 5528 91560 5556
rect 84252 5516 84258 5528
rect 91554 5516 91560 5528
rect 91612 5516 91618 5568
rect 247586 5516 247592 5568
rect 247644 5556 247650 5568
rect 248414 5556 248420 5568
rect 247644 5528 248420 5556
rect 247644 5516 247650 5528
rect 248414 5516 248420 5528
rect 248472 5516 248478 5568
rect 142246 5312 142252 5364
rect 142304 5352 142310 5364
rect 214466 5352 214472 5364
rect 142304 5324 214472 5352
rect 142304 5312 142310 5324
rect 214466 5312 214472 5324
rect 214524 5312 214530 5364
rect 142154 5244 142160 5296
rect 142212 5284 142218 5296
rect 218146 5284 218152 5296
rect 142212 5256 218152 5284
rect 142212 5244 142218 5256
rect 218146 5244 218152 5256
rect 218204 5244 218210 5296
rect 258074 5244 258080 5296
rect 258132 5284 258138 5296
rect 290182 5284 290188 5296
rect 258132 5256 290188 5284
rect 258132 5244 258138 5256
rect 290182 5244 290188 5256
rect 290240 5244 290246 5296
rect 208486 5176 208492 5228
rect 208544 5216 208550 5228
rect 515950 5216 515956 5228
rect 208544 5188 515956 5216
rect 208544 5176 208550 5188
rect 515950 5176 515956 5188
rect 516008 5176 516014 5228
rect 208394 5108 208400 5160
rect 208452 5148 208458 5160
rect 519538 5148 519544 5160
rect 208452 5120 519544 5148
rect 208452 5108 208458 5120
rect 519538 5108 519544 5120
rect 519596 5108 519602 5160
rect 56686 5040 56692 5092
rect 56744 5080 56750 5092
rect 79686 5080 79692 5092
rect 56744 5052 79692 5080
rect 56744 5040 56750 5052
rect 79686 5040 79692 5052
rect 79744 5040 79750 5092
rect 136726 5040 136732 5092
rect 136784 5080 136790 5092
rect 189718 5080 189724 5092
rect 136784 5052 189724 5080
rect 136784 5040 136790 5052
rect 189718 5040 189724 5052
rect 189776 5040 189782 5092
rect 209774 5040 209780 5092
rect 209832 5080 209838 5092
rect 526622 5080 526628 5092
rect 209832 5052 526628 5080
rect 209832 5040 209838 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 56594 4972 56600 5024
rect 56652 5012 56658 5024
rect 83274 5012 83280 5024
rect 56652 4984 83280 5012
rect 56652 4972 56658 4984
rect 83274 4972 83280 4984
rect 83332 4972 83338 5024
rect 136634 4972 136640 5024
rect 136692 5012 136698 5024
rect 193306 5012 193312 5024
rect 136692 4984 193312 5012
rect 136692 4972 136698 4984
rect 193306 4972 193312 4984
rect 193364 4972 193370 5024
rect 211154 4972 211160 5024
rect 211212 5012 211218 5024
rect 530118 5012 530124 5024
rect 211212 4984 530124 5012
rect 211212 4972 211218 4984
rect 530118 4972 530124 4984
rect 530176 4972 530182 5024
rect 57974 4904 57980 4956
rect 58032 4944 58038 4956
rect 86862 4944 86868 4956
rect 58032 4916 86868 4944
rect 58032 4904 58038 4916
rect 86862 4904 86868 4916
rect 86920 4904 86926 4956
rect 138014 4904 138020 4956
rect 138072 4944 138078 4956
rect 196802 4944 196808 4956
rect 138072 4916 196808 4944
rect 138072 4904 138078 4916
rect 196802 4904 196808 4916
rect 196860 4904 196866 4956
rect 212626 4904 212632 4956
rect 212684 4944 212690 4956
rect 533706 4944 533712 4956
rect 212684 4916 533712 4944
rect 212684 4904 212690 4916
rect 533706 4904 533712 4916
rect 533764 4904 533770 4956
rect 62206 4836 62212 4888
rect 62264 4876 62270 4888
rect 104526 4876 104532 4888
rect 62264 4848 104532 4876
rect 62264 4836 62270 4848
rect 104526 4836 104532 4848
rect 104584 4836 104590 4888
rect 138106 4836 138112 4888
rect 138164 4876 138170 4888
rect 200298 4876 200304 4888
rect 138164 4848 200304 4876
rect 138164 4836 138170 4848
rect 200298 4836 200304 4848
rect 200356 4836 200362 4888
rect 212534 4836 212540 4888
rect 212592 4876 212598 4888
rect 537202 4876 537208 4888
rect 212592 4848 537208 4876
rect 212592 4836 212598 4848
rect 537202 4836 537208 4848
rect 537260 4836 537266 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 39298 4808 39304 4820
rect 624 4780 39304 4808
rect 624 4768 630 4780
rect 39298 4768 39304 4780
rect 39356 4768 39362 4820
rect 52454 4768 52460 4820
rect 52512 4808 52518 4820
rect 62022 4808 62028 4820
rect 52512 4780 62028 4808
rect 52512 4768 52518 4780
rect 62022 4768 62028 4780
rect 62080 4768 62086 4820
rect 62114 4768 62120 4820
rect 62172 4808 62178 4820
rect 108114 4808 108120 4820
rect 62172 4780 108120 4808
rect 62172 4768 62178 4780
rect 108114 4768 108120 4780
rect 108172 4768 108178 4820
rect 140774 4768 140780 4820
rect 140832 4808 140838 4820
rect 210970 4808 210976 4820
rect 140832 4780 210976 4808
rect 140832 4768 140838 4780
rect 210970 4768 210976 4780
rect 211028 4768 211034 4820
rect 540790 4808 540796 4820
rect 222166 4780 540796 4808
rect 213914 4700 213920 4752
rect 213972 4740 213978 4752
rect 222166 4740 222194 4780
rect 540790 4768 540796 4780
rect 540848 4768 540854 4820
rect 213972 4712 222194 4740
rect 213972 4700 213978 4712
rect 40678 4564 40684 4616
rect 40736 4604 40742 4616
rect 47578 4604 47584 4616
rect 40736 4576 47584 4604
rect 40736 4564 40742 4576
rect 47578 4564 47584 4576
rect 47636 4564 47642 4616
rect 251266 4496 251272 4548
rect 251324 4536 251330 4548
rect 258258 4536 258264 4548
rect 251324 4508 258264 4536
rect 251324 4496 251330 4508
rect 258258 4496 258264 4508
rect 258316 4496 258322 4548
rect 82814 4292 82820 4344
rect 82872 4332 82878 4344
rect 84470 4332 84476 4344
rect 82872 4304 84476 4332
rect 82872 4292 82878 4304
rect 84470 4292 84476 4304
rect 84528 4292 84534 4344
rect 49694 4224 49700 4276
rect 49752 4264 49758 4276
rect 51350 4264 51356 4276
rect 49752 4236 51356 4264
rect 49752 4224 49758 4236
rect 51350 4224 51356 4236
rect 51408 4224 51414 4276
rect 47854 4156 47860 4208
rect 47912 4196 47918 4208
rect 49786 4196 49792 4208
rect 47912 4168 49792 4196
rect 47912 4156 47918 4168
rect 49786 4156 49792 4168
rect 49844 4156 49850 4208
rect 51074 4156 51080 4208
rect 51132 4196 51138 4208
rect 54938 4196 54944 4208
rect 51132 4168 54944 4196
rect 51132 4156 51138 4168
rect 54938 4156 54944 4168
rect 54996 4156 55002 4208
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 17218 4128 17224 4140
rect 14792 4100 17224 4128
rect 14792 4088 14798 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 97994 4128 98000 4140
rect 43128 4100 98000 4128
rect 43128 4088 43134 4100
rect 97994 4088 98000 4100
rect 98052 4088 98058 4140
rect 323302 4088 323308 4140
rect 323360 4128 323366 4140
rect 364518 4128 364524 4140
rect 323360 4100 364524 4128
rect 323360 4088 323366 4100
rect 364518 4088 364524 4100
rect 364576 4088 364582 4140
rect 389174 4088 389180 4140
rect 389232 4128 389238 4140
rect 436738 4128 436744 4140
rect 389232 4100 436744 4128
rect 389232 4088 389238 4100
rect 436738 4088 436744 4100
rect 436796 4088 436802 4140
rect 39574 4020 39580 4072
rect 39632 4060 39638 4072
rect 98086 4060 98092 4072
rect 39632 4032 98092 4060
rect 39632 4020 39638 4032
rect 98086 4020 98092 4032
rect 98144 4020 98150 4072
rect 319714 4020 319720 4072
rect 319772 4060 319778 4072
rect 364426 4060 364432 4072
rect 319772 4032 364432 4060
rect 319772 4020 319778 4032
rect 364426 4020 364432 4032
rect 364484 4020 364490 4072
rect 390554 4020 390560 4072
rect 390612 4060 390618 4072
rect 440234 4060 440240 4072
rect 390612 4032 440240 4060
rect 390612 4020 390618 4032
rect 440234 4020 440240 4032
rect 440292 4020 440298 4072
rect 35986 3952 35992 4004
rect 36044 3992 36050 4004
rect 96706 3992 96712 4004
rect 36044 3964 96712 3992
rect 36044 3952 36050 3964
rect 96706 3952 96712 3964
rect 96764 3952 96770 4004
rect 316218 3952 316224 4004
rect 316276 3992 316282 4004
rect 362954 3992 362960 4004
rect 316276 3964 362960 3992
rect 316276 3952 316282 3964
rect 362954 3952 362960 3964
rect 363012 3952 363018 4004
rect 391934 3952 391940 4004
rect 391992 3992 391998 4004
rect 443822 3992 443828 4004
rect 391992 3964 443828 3992
rect 391992 3952 391998 3964
rect 443822 3952 443828 3964
rect 443880 3952 443886 4004
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 96614 3924 96620 3936
rect 32456 3896 96620 3924
rect 32456 3884 32462 3896
rect 96614 3884 96620 3896
rect 96672 3884 96678 3936
rect 121638 3884 121644 3936
rect 121696 3924 121702 3936
rect 125870 3924 125876 3936
rect 121696 3896 125876 3924
rect 121696 3884 121702 3896
rect 125870 3884 125876 3896
rect 125928 3884 125934 3936
rect 312630 3884 312636 3936
rect 312688 3924 312694 3936
rect 363046 3924 363052 3936
rect 312688 3896 363052 3924
rect 312688 3884 312694 3896
rect 363046 3884 363052 3896
rect 363104 3884 363110 3936
rect 385034 3884 385040 3936
rect 385092 3924 385098 3936
rect 392026 3924 392032 3936
rect 385092 3896 392032 3924
rect 385092 3884 385098 3896
rect 392026 3884 392032 3896
rect 392084 3884 392090 3936
rect 393314 3884 393320 3936
rect 393372 3924 393378 3936
rect 450906 3924 450912 3936
rect 393372 3896 450912 3924
rect 393372 3884 393378 3896
rect 450906 3884 450912 3896
rect 450964 3884 450970 3936
rect 28902 3816 28908 3868
rect 28960 3856 28966 3868
rect 95326 3856 95332 3868
rect 28960 3828 95332 3856
rect 28960 3816 28966 3828
rect 95326 3816 95332 3828
rect 95384 3816 95390 3868
rect 103330 3816 103336 3868
rect 103388 3856 103394 3868
rect 111886 3856 111892 3868
rect 103388 3828 111892 3856
rect 103388 3816 103394 3828
rect 111886 3816 111892 3828
rect 111944 3816 111950 3868
rect 120166 3856 120172 3868
rect 113146 3828 120172 3856
rect 24210 3748 24216 3800
rect 24268 3788 24274 3800
rect 95234 3788 95240 3800
rect 24268 3760 95240 3788
rect 24268 3748 24274 3760
rect 95234 3748 95240 3760
rect 95292 3748 95298 3800
rect 99834 3748 99840 3800
rect 99892 3788 99898 3800
rect 111794 3788 111800 3800
rect 99892 3760 111800 3788
rect 99892 3748 99898 3760
rect 111794 3748 111800 3760
rect 111852 3748 111858 3800
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 94038 3720 94044 3732
rect 19484 3692 94044 3720
rect 19484 3680 19490 3692
rect 94038 3680 94044 3692
rect 94096 3680 94102 3732
rect 96246 3680 96252 3732
rect 96304 3720 96310 3732
rect 110598 3720 110604 3732
rect 96304 3692 110604 3720
rect 96304 3680 96310 3692
rect 110598 3680 110604 3692
rect 110656 3680 110662 3732
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 113146 3652 113174 3828
rect 120166 3816 120172 3828
rect 120224 3816 120230 3868
rect 168374 3816 168380 3868
rect 168432 3856 168438 3868
rect 169570 3856 169576 3868
rect 168432 3828 169576 3856
rect 168432 3816 168438 3828
rect 169570 3816 169576 3828
rect 169628 3816 169634 3868
rect 176746 3816 176752 3868
rect 176804 3856 176810 3868
rect 177850 3856 177856 3868
rect 176804 3828 177856 3856
rect 176804 3816 176810 3828
rect 177850 3816 177856 3828
rect 177908 3816 177914 3868
rect 251174 3816 251180 3868
rect 251232 3856 251238 3868
rect 252370 3856 252376 3868
rect 251232 3828 252376 3856
rect 251232 3816 251238 3828
rect 252370 3816 252376 3828
rect 252428 3816 252434 3868
rect 291378 3816 291384 3868
rect 291436 3856 291442 3868
rect 294598 3856 294604 3868
rect 291436 3828 294604 3856
rect 291436 3816 291442 3828
rect 294598 3816 294604 3828
rect 294656 3816 294662 3868
rect 309042 3816 309048 3868
rect 309100 3856 309106 3868
rect 361666 3856 361672 3868
rect 309100 3828 361672 3856
rect 309100 3816 309106 3828
rect 361666 3816 361672 3828
rect 361724 3816 361730 3868
rect 362310 3816 362316 3868
rect 362368 3856 362374 3868
rect 373994 3856 374000 3868
rect 362368 3828 374000 3856
rect 362368 3816 362374 3828
rect 373994 3816 374000 3828
rect 374052 3816 374058 3868
rect 379514 3816 379520 3868
rect 379572 3856 379578 3868
rect 387150 3856 387156 3868
rect 379572 3828 387156 3856
rect 379572 3816 379578 3828
rect 387150 3816 387156 3828
rect 387208 3816 387214 3868
rect 394694 3816 394700 3868
rect 394752 3856 394758 3868
rect 458082 3856 458088 3868
rect 394752 3828 458088 3856
rect 394752 3816 394758 3828
rect 458082 3816 458088 3828
rect 458140 3816 458146 3868
rect 160094 3748 160100 3800
rect 160152 3788 160158 3800
rect 328546 3788 328552 3800
rect 160152 3760 328552 3788
rect 160152 3748 160158 3760
rect 328546 3748 328552 3760
rect 328604 3748 328610 3800
rect 348050 3748 348056 3800
rect 348108 3788 348114 3800
rect 369946 3788 369952 3800
rect 348108 3760 369952 3788
rect 348108 3748 348114 3760
rect 369946 3748 369952 3760
rect 370004 3748 370010 3800
rect 379606 3748 379612 3800
rect 379664 3788 379670 3800
rect 390554 3788 390560 3800
rect 379664 3760 390560 3788
rect 379664 3748 379670 3760
rect 390554 3748 390560 3760
rect 390612 3748 390618 3800
rect 396074 3748 396080 3800
rect 396132 3788 396138 3800
rect 465166 3788 465172 3800
rect 396132 3760 465172 3788
rect 396132 3748 396138 3760
rect 465166 3748 465172 3760
rect 465224 3748 465230 3800
rect 124306 3680 124312 3732
rect 124364 3720 124370 3732
rect 132954 3720 132960 3732
rect 124364 3692 132960 3720
rect 124364 3680 124370 3692
rect 132954 3680 132960 3692
rect 133012 3680 133018 3732
rect 135254 3680 135260 3732
rect 135312 3720 135318 3732
rect 140038 3720 140044 3732
rect 135312 3692 140044 3720
rect 135312 3680 135318 3692
rect 140038 3680 140044 3692
rect 140096 3680 140102 3732
rect 156598 3680 156604 3732
rect 156656 3720 156662 3732
rect 328454 3720 328460 3732
rect 156656 3692 328460 3720
rect 156656 3680 156662 3692
rect 328454 3680 328460 3692
rect 328512 3680 328518 3732
rect 344554 3680 344560 3732
rect 344612 3720 344618 3732
rect 369854 3720 369860 3732
rect 344612 3692 369860 3720
rect 344612 3680 344618 3692
rect 369854 3680 369860 3692
rect 369912 3680 369918 3732
rect 372890 3680 372896 3732
rect 372948 3720 372954 3732
rect 375558 3720 375564 3732
rect 372948 3692 375564 3720
rect 372948 3680 372954 3692
rect 375558 3680 375564 3692
rect 375616 3680 375622 3732
rect 380894 3680 380900 3732
rect 380952 3720 380958 3732
rect 394234 3720 394240 3732
rect 380952 3692 394240 3720
rect 380952 3680 380958 3692
rect 394234 3680 394240 3692
rect 394292 3680 394298 3732
rect 397454 3680 397460 3732
rect 397512 3720 397518 3732
rect 472250 3720 472256 3732
rect 397512 3692 472256 3720
rect 397512 3680 397518 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 118970 3652 118976 3664
rect 25372 3624 113174 3652
rect 115400 3624 118976 3652
rect 25372 3612 25378 3624
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 15838 3584 15844 3596
rect 10008 3556 15844 3584
rect 10008 3544 10014 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 115400 3584 115428 3624
rect 118970 3612 118976 3624
rect 119028 3612 119034 3664
rect 124214 3612 124220 3664
rect 124272 3652 124278 3664
rect 136450 3652 136456 3664
rect 124272 3624 136456 3652
rect 124272 3612 124278 3624
rect 136450 3612 136456 3624
rect 136508 3612 136514 3664
rect 153010 3612 153016 3664
rect 153068 3652 153074 3664
rect 327166 3652 327172 3664
rect 153068 3624 327172 3652
rect 153068 3612 153074 3624
rect 327166 3612 327172 3624
rect 327224 3612 327230 3664
rect 337470 3612 337476 3664
rect 337528 3652 337534 3664
rect 368566 3652 368572 3664
rect 337528 3624 368572 3652
rect 337528 3612 337534 3624
rect 368566 3612 368572 3624
rect 368624 3612 368630 3664
rect 385126 3612 385132 3664
rect 385184 3652 385190 3664
rect 407022 3652 407028 3664
rect 385184 3624 407028 3652
rect 385184 3612 385190 3624
rect 407022 3612 407028 3624
rect 407080 3612 407086 3664
rect 407206 3612 407212 3664
rect 407264 3652 407270 3664
rect 408402 3652 408408 3664
rect 407264 3624 408408 3652
rect 407264 3612 407270 3624
rect 408402 3612 408408 3624
rect 408460 3612 408466 3664
rect 415394 3652 415400 3664
rect 412606 3624 415400 3652
rect 118694 3584 118700 3596
rect 20680 3556 115428 3584
rect 116044 3556 118700 3584
rect 20680 3544 20686 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4798 3516 4804 3528
rect 2924 3488 4804 3516
rect 2924 3476 2930 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 116044 3516 116072 3556
rect 118694 3544 118700 3556
rect 118752 3544 118758 3596
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 147122 3584 147128 3596
rect 127032 3556 147128 3584
rect 127032 3544 127038 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 149514 3544 149520 3596
rect 149572 3584 149578 3596
rect 327258 3584 327264 3596
rect 149572 3556 327264 3584
rect 149572 3544 149578 3556
rect 327258 3544 327264 3556
rect 327316 3544 327322 3596
rect 333882 3544 333888 3596
rect 333940 3584 333946 3596
rect 367094 3584 367100 3596
rect 333940 3556 367100 3584
rect 333940 3544 333946 3556
rect 367094 3544 367100 3556
rect 367152 3544 367158 3596
rect 386414 3544 386420 3596
rect 386472 3584 386478 3596
rect 386472 3556 391980 3584
rect 386472 3544 386478 3556
rect 15988 3488 116072 3516
rect 15988 3476 15994 3488
rect 116578 3476 116584 3528
rect 116636 3516 116642 3528
rect 117590 3516 117596 3528
rect 116636 3488 117596 3516
rect 116636 3476 116642 3488
rect 117590 3476 117596 3488
rect 117648 3476 117654 3528
rect 128170 3476 128176 3528
rect 128228 3516 128234 3528
rect 129090 3516 129096 3528
rect 128228 3488 129096 3516
rect 128228 3476 128234 3488
rect 129090 3476 129096 3488
rect 129148 3476 129154 3528
rect 143534 3516 143540 3528
rect 129200 3488 143540 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 10318 3448 10324 3460
rect 6512 3420 10324 3448
rect 6512 3408 6518 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 117314 3448 117320 3460
rect 11204 3420 117320 3448
rect 11204 3408 11210 3420
rect 117314 3408 117320 3420
rect 117372 3408 117378 3460
rect 125594 3408 125600 3460
rect 125652 3448 125658 3460
rect 129200 3448 129228 3488
rect 143534 3476 143540 3488
rect 143592 3476 143598 3528
rect 145926 3476 145932 3528
rect 145984 3516 145990 3528
rect 325694 3516 325700 3528
rect 145984 3488 325700 3516
rect 145984 3476 145990 3488
rect 325694 3476 325700 3488
rect 325752 3476 325758 3528
rect 330386 3476 330392 3528
rect 330444 3516 330450 3528
rect 365714 3516 365720 3528
rect 330444 3488 365720 3516
rect 330444 3476 330450 3488
rect 365714 3476 365720 3488
rect 365772 3476 365778 3528
rect 390646 3476 390652 3528
rect 390704 3516 390710 3528
rect 391842 3516 391848 3528
rect 390704 3488 391848 3516
rect 390704 3476 390710 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 391952 3516 391980 3556
rect 392026 3544 392032 3596
rect 392084 3584 392090 3596
rect 412606 3584 412634 3624
rect 415394 3612 415400 3624
rect 415452 3612 415458 3664
rect 423582 3612 423588 3664
rect 423640 3652 423646 3664
rect 582190 3652 582196 3664
rect 423640 3624 582196 3652
rect 423640 3612 423646 3624
rect 582190 3612 582196 3624
rect 582248 3612 582254 3664
rect 418982 3584 418988 3596
rect 392084 3556 412634 3584
rect 415412 3556 418988 3584
rect 392084 3544 392090 3556
rect 415412 3516 415440 3556
rect 418982 3544 418988 3556
rect 419040 3544 419046 3596
rect 420914 3544 420920 3596
rect 420972 3584 420978 3596
rect 578602 3584 578608 3596
rect 420972 3556 578608 3584
rect 420972 3544 420978 3556
rect 578602 3544 578608 3556
rect 578660 3544 578666 3596
rect 391952 3488 415440 3516
rect 415486 3476 415492 3528
rect 415544 3516 415550 3528
rect 416682 3516 416688 3528
rect 415544 3488 416688 3516
rect 415544 3476 415550 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 422386 3476 422392 3528
rect 422444 3516 422450 3528
rect 580994 3516 581000 3528
rect 422444 3488 581000 3516
rect 422444 3476 422450 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 140038 3448 140044 3460
rect 125652 3420 129228 3448
rect 132466 3420 140044 3448
rect 125652 3408 125658 3420
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 99374 3380 99380 3392
rect 46716 3352 99380 3380
rect 46716 3340 46722 3352
rect 99374 3340 99380 3352
rect 99432 3340 99438 3392
rect 125686 3340 125692 3392
rect 125744 3380 125750 3392
rect 132466 3380 132494 3420
rect 140038 3408 140044 3420
rect 140096 3408 140102 3460
rect 142430 3408 142436 3460
rect 142488 3448 142494 3460
rect 325786 3448 325792 3460
rect 142488 3420 325792 3448
rect 142488 3408 142494 3420
rect 325786 3408 325792 3420
rect 325844 3408 325850 3460
rect 326798 3408 326804 3460
rect 326856 3448 326862 3460
rect 326856 3420 365116 3448
rect 326856 3408 326862 3420
rect 125744 3352 132494 3380
rect 125744 3340 125750 3352
rect 193214 3340 193220 3392
rect 193272 3380 193278 3392
rect 194410 3380 194416 3392
rect 193272 3352 194416 3380
rect 193272 3340 193278 3352
rect 194410 3340 194416 3352
rect 194468 3340 194474 3392
rect 287790 3340 287796 3392
rect 287848 3380 287854 3392
rect 291838 3380 291844 3392
rect 287848 3352 291844 3380
rect 287848 3340 287854 3352
rect 291838 3340 291844 3352
rect 291896 3340 291902 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 351638 3340 351644 3392
rect 351696 3380 351702 3392
rect 365088 3380 365116 3420
rect 365806 3408 365812 3460
rect 365864 3448 365870 3460
rect 374178 3448 374184 3460
rect 365864 3420 374184 3448
rect 365864 3408 365870 3420
rect 374178 3408 374184 3420
rect 374236 3408 374242 3460
rect 386506 3408 386512 3460
rect 386564 3448 386570 3460
rect 422570 3448 422576 3460
rect 386564 3420 422576 3448
rect 386564 3408 386570 3420
rect 422570 3408 422576 3420
rect 422628 3408 422634 3460
rect 423674 3408 423680 3460
rect 423732 3448 423738 3460
rect 583386 3448 583392 3460
rect 423732 3420 583392 3448
rect 423732 3408 423738 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 365898 3380 365904 3392
rect 351696 3352 365024 3380
rect 365088 3352 365904 3380
rect 351696 3340 351702 3352
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 109034 3312 109040 3324
rect 89220 3284 109040 3312
rect 89220 3272 89226 3284
rect 109034 3272 109040 3284
rect 109092 3272 109098 3324
rect 116026 3272 116032 3324
rect 116084 3312 116090 3324
rect 124674 3312 124680 3324
rect 116084 3284 124680 3312
rect 116084 3272 116090 3284
rect 124674 3272 124680 3284
rect 124732 3272 124738 3324
rect 355226 3272 355232 3324
rect 355284 3312 355290 3324
rect 364996 3312 365024 3352
rect 365898 3340 365904 3352
rect 365956 3340 365962 3392
rect 389266 3340 389272 3392
rect 389324 3380 389330 3392
rect 433242 3380 433248 3392
rect 389324 3352 433248 3380
rect 389324 3340 389330 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 523034 3340 523040 3392
rect 523092 3380 523098 3392
rect 523862 3380 523868 3392
rect 523092 3352 523868 3380
rect 523092 3340 523098 3352
rect 523862 3340 523868 3352
rect 523920 3340 523926 3392
rect 547874 3340 547880 3392
rect 547932 3380 547938 3392
rect 548702 3380 548708 3392
rect 547932 3352 548708 3380
rect 547932 3340 547938 3352
rect 548702 3340 548708 3352
rect 548760 3340 548766 3392
rect 564434 3340 564440 3392
rect 564492 3380 564498 3392
rect 565262 3380 565268 3392
rect 564492 3352 565268 3380
rect 564492 3340 564498 3352
rect 565262 3340 565268 3352
rect 565320 3340 565326 3392
rect 371234 3312 371240 3324
rect 355284 3284 364932 3312
rect 364996 3284 371240 3312
rect 355284 3272 355290 3284
rect 92750 3204 92756 3256
rect 92808 3244 92814 3256
rect 109126 3244 109132 3256
rect 92808 3216 109132 3244
rect 92808 3204 92814 3216
rect 109126 3204 109132 3216
rect 109184 3204 109190 3256
rect 122926 3204 122932 3256
rect 122984 3244 122990 3256
rect 129366 3244 129372 3256
rect 122984 3216 129372 3244
rect 122984 3204 122990 3216
rect 129366 3204 129372 3216
rect 129424 3204 129430 3256
rect 364904 3244 364932 3284
rect 371234 3272 371240 3284
rect 371292 3272 371298 3324
rect 376938 3272 376944 3324
rect 376996 3312 377002 3324
rect 379974 3312 379980 3324
rect 376996 3284 379980 3312
rect 376996 3272 377002 3284
rect 379974 3272 379980 3284
rect 380032 3272 380038 3324
rect 387886 3272 387892 3324
rect 387944 3312 387950 3324
rect 429654 3312 429660 3324
rect 387944 3284 429660 3312
rect 387944 3272 387950 3284
rect 429654 3272 429660 3284
rect 429712 3272 429718 3324
rect 371326 3244 371332 3256
rect 364904 3216 371332 3244
rect 371326 3204 371332 3216
rect 371384 3204 371390 3256
rect 387794 3204 387800 3256
rect 387852 3244 387858 3256
rect 426158 3244 426164 3256
rect 387852 3216 426164 3244
rect 387852 3204 387858 3216
rect 426158 3204 426164 3216
rect 426216 3204 426222 3256
rect 369394 3136 369400 3188
rect 369452 3176 369458 3188
rect 375466 3176 375472 3188
rect 369452 3148 375472 3176
rect 369452 3136 369458 3148
rect 375466 3136 375472 3148
rect 375524 3136 375530 3188
rect 407022 3136 407028 3188
rect 407080 3176 407086 3188
rect 411898 3176 411904 3188
rect 407080 3148 411904 3176
rect 407080 3136 407086 3148
rect 411898 3136 411904 3148
rect 411956 3136 411962 3188
rect 115934 3068 115940 3120
rect 115992 3108 115998 3120
rect 121086 3108 121092 3120
rect 115992 3080 121092 3108
rect 115992 3068 115998 3080
rect 121086 3068 121092 3080
rect 121144 3068 121150 3120
rect 358722 3068 358728 3120
rect 358780 3108 358786 3120
rect 372614 3108 372620 3120
rect 358780 3080 372620 3108
rect 358780 3068 358786 3080
rect 372614 3068 372620 3080
rect 372672 3068 372678 3120
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 3970 3040 3976 3052
rect 1728 3012 3976 3040
rect 1728 3000 1734 3012
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 378134 2932 378140 2984
rect 378192 2972 378198 2984
rect 383562 2972 383568 2984
rect 378192 2944 383568 2972
rect 378192 2932 378198 2944
rect 383562 2932 383568 2944
rect 383620 2932 383626 2984
rect 301958 2864 301964 2916
rect 302016 2904 302022 2916
rect 307018 2904 307024 2916
rect 302016 2876 307024 2904
rect 302016 2864 302022 2876
rect 307018 2864 307024 2876
rect 307076 2864 307082 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 314660 700952 314712 701004
rect 413652 700952 413704 701004
rect 325700 700884 325752 700936
rect 429844 700884 429896 700936
rect 336740 700816 336792 700868
rect 446128 700816 446180 700868
rect 347872 700748 347924 700800
rect 462320 700748 462372 700800
rect 358820 700680 358872 700732
rect 478512 700680 478564 700732
rect 248420 700612 248472 700664
rect 316316 700612 316368 700664
rect 369860 700612 369912 700664
rect 494796 700612 494848 700664
rect 259460 700544 259512 700596
rect 332508 700544 332560 700596
rect 379520 700544 379572 700596
rect 510988 700544 511040 700596
rect 204260 700476 204312 700528
rect 251456 700476 251508 700528
rect 270500 700476 270552 700528
rect 348792 700476 348844 700528
rect 390560 700476 390612 700528
rect 527180 700476 527232 700528
rect 171140 700408 171192 700460
rect 202788 700408 202840 700460
rect 215300 700408 215352 700460
rect 267648 700408 267700 700460
rect 281540 700408 281592 700460
rect 364984 700408 365036 700460
rect 401600 700408 401652 700460
rect 543464 700408 543516 700460
rect 149060 700340 149112 700392
rect 170312 700340 170364 700392
rect 182180 700340 182232 700392
rect 218980 700340 219032 700392
rect 226340 700340 226392 700392
rect 283840 700340 283892 700392
rect 292580 700340 292632 700392
rect 381176 700340 381228 700392
rect 412640 700340 412692 700392
rect 559656 700340 559708 700392
rect 126980 700272 127032 700324
rect 137836 700272 137888 700324
rect 138020 700272 138072 700324
rect 154120 700272 154172 700324
rect 160100 700272 160152 700324
rect 186504 700272 186556 700324
rect 193220 700272 193272 700324
rect 235172 700272 235224 700324
rect 237380 700272 237432 700324
rect 300124 700272 300176 700324
rect 303620 700272 303672 700324
rect 397460 700272 397512 700324
rect 423680 700272 423732 700324
rect 575848 700272 575900 700324
rect 115940 699660 115992 699712
rect 121644 699660 121696 699712
rect 3424 683748 3476 683800
rect 11704 683748 11756 683800
rect 428464 683136 428516 683188
rect 579620 683136 579672 683188
rect 3516 670964 3568 671016
rect 4804 670964 4856 671016
rect 3516 656888 3568 656940
rect 33784 656888 33836 656940
rect 2872 644444 2924 644496
rect 10324 644444 10376 644496
rect 3516 632068 3568 632120
rect 22744 632068 22796 632120
rect 428556 630640 428608 630692
rect 579620 630640 579672 630692
rect 3332 605820 3384 605872
rect 36544 605820 36596 605872
rect 3332 592016 3384 592068
rect 14464 592016 14516 592068
rect 3332 579640 3384 579692
rect 25504 579640 25556 579692
rect 428648 576852 428700 576904
rect 580172 576852 580224 576904
rect 88340 562980 88392 563032
rect 94596 562980 94648 563032
rect 40040 562436 40092 562488
rect 61660 562436 61712 562488
rect 71780 562436 71832 562488
rect 83648 562436 83700 562488
rect 23480 562368 23532 562420
rect 50620 562368 50672 562420
rect 6920 562300 6972 562352
rect 40408 562300 40460 562352
rect 56600 562300 56652 562352
rect 72700 562300 72752 562352
rect 3148 553528 3200 553580
rect 6184 553528 6236 553580
rect 490564 550604 490616 550656
rect 580172 550604 580224 550656
rect 11704 545028 11756 545080
rect 37832 545028 37884 545080
rect 428740 545028 428792 545080
rect 580264 545028 580316 545080
rect 22744 541628 22796 541680
rect 37924 541628 37976 541680
rect 3056 539588 3108 539640
rect 22744 539588 22796 539640
rect 4804 536732 4856 536784
rect 37556 536732 37608 536784
rect 2964 527144 3016 527196
rect 28264 527144 28316 527196
rect 3424 527076 3476 527128
rect 37832 527076 37884 527128
rect 428740 525716 428792 525768
rect 580356 525716 580408 525768
rect 428464 524424 428516 524476
rect 580172 524424 580224 524476
rect 33784 517420 33836 517472
rect 38016 517420 38068 517472
rect 428740 516060 428792 516112
rect 580448 516060 580500 516112
rect 10324 507764 10376 507816
rect 37556 507764 37608 507816
rect 428740 506404 428792 506456
rect 580540 506404 580592 506456
rect 3148 488520 3200 488572
rect 10324 488520 10376 488572
rect 3516 488452 3568 488504
rect 37832 488452 37884 488504
rect 428556 487092 428608 487144
rect 580632 487092 580684 487144
rect 428556 477436 428608 477488
rect 580724 477436 580776 477488
rect 3516 474716 3568 474768
rect 31024 474716 31076 474768
rect 428556 470568 428608 470620
rect 579988 470568 580040 470620
rect 14464 469140 14516 469192
rect 37924 469140 37976 469192
rect 428740 467780 428792 467832
rect 580724 467780 580776 467832
rect 25504 459484 25556 459536
rect 37464 459484 37516 459536
rect 3608 449828 3660 449880
rect 37924 449828 37976 449880
rect 429108 448468 429160 448520
rect 580908 448468 580960 448520
rect 6184 441532 6236 441584
rect 37832 441532 37884 441584
rect 428648 438812 428700 438864
rect 490564 438812 490616 438864
rect 3332 436092 3384 436144
rect 11704 436092 11756 436144
rect 22744 431876 22796 431928
rect 37832 431876 37884 431928
rect 428740 430584 428792 430636
rect 580080 430584 580132 430636
rect 428648 429088 428700 429140
rect 580264 429088 580316 429140
rect 3332 422288 3384 422340
rect 26884 422288 26936 422340
rect 28264 422220 28316 422272
rect 37924 422220 37976 422272
rect 428740 418140 428792 418192
rect 580172 418140 580224 418192
rect 3424 412564 3476 412616
rect 37648 412564 37700 412616
rect 428832 409776 428884 409828
rect 580356 409776 580408 409828
rect 3700 402908 3752 402960
rect 37556 402908 37608 402960
rect 428464 400120 428516 400172
rect 580448 400120 580500 400172
rect 10324 393252 10376 393304
rect 37740 393252 37792 393304
rect 428464 390464 428516 390516
rect 580540 390464 580592 390516
rect 3332 383664 3384 383716
rect 24124 383664 24176 383716
rect 31024 383596 31076 383648
rect 37464 383596 37516 383648
rect 3516 373940 3568 373992
rect 37924 373940 37976 373992
rect 3148 371288 3200 371340
rect 6184 371288 6236 371340
rect 428832 371152 428884 371204
rect 580632 371152 580684 371204
rect 428464 364352 428516 364404
rect 579804 364352 579856 364404
rect 3792 364284 3844 364336
rect 37464 364284 37516 364336
rect 428556 361496 428608 361548
rect 580724 361496 580776 361548
rect 11704 354628 11756 354680
rect 37556 354628 37608 354680
rect 26884 344972 26936 345024
rect 37648 344972 37700 345024
rect 3424 336676 3476 336728
rect 37832 336676 37884 336728
rect 428556 332528 428608 332580
rect 580264 332528 580316 332580
rect 2780 331576 2832 331628
rect 4804 331576 4856 331628
rect 3608 327020 3660 327072
rect 37556 327020 37608 327072
rect 428556 324300 428608 324352
rect 579620 324300 579672 324352
rect 428832 322872 428884 322924
rect 580356 322872 580408 322924
rect 24124 317364 24176 317416
rect 37924 317364 37976 317416
rect 428740 313216 428792 313268
rect 580448 313216 580500 313268
rect 428648 311856 428700 311908
rect 580172 311856 580224 311908
rect 6184 307708 6236 307760
rect 37372 307708 37424 307760
rect 3516 298052 3568 298104
rect 37556 298052 37608 298104
rect 428464 292476 428516 292528
rect 580540 292476 580592 292528
rect 3700 288328 3752 288380
rect 37740 288328 37792 288380
rect 429016 282820 429068 282872
rect 580632 282820 580684 282872
rect 4804 278672 4856 278724
rect 37740 278672 37792 278724
rect 428464 271872 428516 271924
rect 579620 271872 579672 271924
rect 3424 269016 3476 269068
rect 37924 269016 37976 269068
rect 3608 259360 3660 259412
rect 37372 259360 37424 259412
rect 428556 258068 428608 258120
rect 579620 258068 579672 258120
rect 428924 253852 428976 253904
rect 580264 253852 580316 253904
rect 3516 249704 3568 249756
rect 37924 249704 37976 249756
rect 428740 244264 428792 244316
rect 579804 244264 579856 244316
rect 428648 244196 428700 244248
rect 580356 244196 580408 244248
rect 3700 240048 3752 240100
rect 37372 240048 37424 240100
rect 428464 231820 428516 231872
rect 580172 231820 580224 231872
rect 3424 231752 3476 231804
rect 37648 231752 37700 231804
rect 3608 222096 3660 222148
rect 37740 222096 37792 222148
rect 428556 218016 428608 218068
rect 580172 218016 580224 218068
rect 3516 212440 3568 212492
rect 37832 212440 37884 212492
rect 428648 205640 428700 205692
rect 580172 205640 580224 205692
rect 3424 202784 3476 202836
rect 37740 202784 37792 202836
rect 3608 193128 3660 193180
rect 37740 193128 37792 193180
rect 428464 191836 428516 191888
rect 580172 191836 580224 191888
rect 3516 183472 3568 183524
rect 37924 183472 37976 183524
rect 428556 178032 428608 178084
rect 580172 178032 580224 178084
rect 3424 173816 3476 173868
rect 37740 173816 37792 173868
rect 428464 165588 428516 165640
rect 580172 165588 580224 165640
rect 3516 164160 3568 164212
rect 37924 164160 37976 164212
rect 3424 154504 3476 154556
rect 37648 154504 37700 154556
rect 429108 151784 429160 151836
rect 579988 151784 580040 151836
rect 3332 144848 3384 144900
rect 37924 144848 37976 144900
rect 428832 137980 428884 138032
rect 580172 137980 580224 138032
rect 3424 136552 3476 136604
rect 37556 136552 37608 136604
rect 428924 126896 428976 126948
rect 580172 126896 580224 126948
rect 3424 124108 3476 124160
rect 37740 124108 37792 124160
rect 428464 113092 428516 113144
rect 579804 113092 579856 113144
rect 3424 111732 3476 111784
rect 37924 111732 37976 111784
rect 428464 100648 428516 100700
rect 580172 100648 580224 100700
rect 3424 97928 3476 97980
rect 37924 97928 37976 97980
rect 428556 86912 428608 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 38016 85484 38068 85536
rect 428464 73108 428516 73160
rect 580172 73108 580224 73160
rect 3424 71680 3476 71732
rect 37924 71680 37976 71732
rect 428556 60664 428608 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 38016 59304 38068 59356
rect 428464 46860 428516 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 37924 45500 37976 45552
rect 212540 39516 212592 39568
rect 212908 39516 212960 39568
rect 72424 38564 72476 38616
rect 73988 38564 74040 38616
rect 194048 38428 194100 38480
rect 195244 38428 195296 38480
rect 297088 38428 297140 38480
rect 312544 38428 312596 38480
rect 55864 38360 55916 38412
rect 58624 38360 58676 38412
rect 207296 38360 207348 38412
rect 209044 38360 209096 38412
rect 311808 38360 311860 38412
rect 349804 38360 349856 38412
rect 47584 38292 47636 38344
rect 48320 38292 48372 38344
rect 282184 38292 282236 38344
rect 324596 38292 324648 38344
rect 324964 38292 325016 38344
rect 356612 38292 356664 38344
rect 411812 38292 411864 38344
rect 425704 38292 425756 38344
rect 46204 38224 46256 38276
rect 48964 38224 49016 38276
rect 185400 38224 185452 38276
rect 188344 38224 188396 38276
rect 203432 38224 203484 38276
rect 224132 38224 224184 38276
rect 286324 38224 286376 38276
rect 330024 38224 330076 38276
rect 330576 38224 330628 38276
rect 348792 38224 348844 38276
rect 375380 38224 375432 38276
rect 376852 38224 376904 38276
rect 393044 38224 393096 38276
rect 447140 38224 447192 38276
rect 75920 38156 75972 38208
rect 77300 38156 77352 38208
rect 163596 38156 163648 38208
rect 170404 38156 170456 38208
rect 171324 38156 171376 38208
rect 172704 38156 172756 38208
rect 181536 38156 181588 38208
rect 218704 38156 218756 38208
rect 226616 38156 226668 38208
rect 244280 38156 244332 38208
rect 277216 38156 277268 38208
rect 307116 38156 307168 38208
rect 322020 38156 322072 38208
rect 414664 38156 414716 38208
rect 415676 38156 415728 38208
rect 436744 38156 436796 38208
rect 66812 38088 66864 38140
rect 68928 38088 68980 38140
rect 169668 38088 169720 38140
rect 200764 38088 200816 38140
rect 215852 38088 215904 38140
rect 342904 38088 342956 38140
rect 394608 38088 394660 38140
rect 454040 38088 454092 38140
rect 59728 38020 59780 38072
rect 69664 38020 69716 38072
rect 84752 38020 84804 38072
rect 86960 38020 87012 38072
rect 91008 38020 91060 38072
rect 93124 38020 93176 38072
rect 98000 38020 98052 38072
rect 99012 38020 99064 38072
rect 101404 38020 101456 38072
rect 102140 38020 102192 38072
rect 39304 37952 39356 38004
rect 40500 37952 40552 38004
rect 41328 37952 41380 38004
rect 41972 37952 42024 38004
rect 44180 37952 44232 38004
rect 45100 37952 45152 38004
rect 49700 37952 49752 38004
rect 50620 37952 50672 38004
rect 52460 37952 52512 38004
rect 52920 37952 52972 38004
rect 56600 37952 56652 38004
rect 57612 37952 57664 38004
rect 62120 37952 62172 38004
rect 63132 37952 63184 38004
rect 64880 37952 64932 38004
rect 65432 37952 65484 38004
rect 70400 37952 70452 38004
rect 70860 37952 70912 38004
rect 71044 37952 71096 38004
rect 73252 37952 73304 38004
rect 74540 37952 74592 38004
rect 75552 37952 75604 38004
rect 80060 37952 80112 38004
rect 80980 37952 81032 38004
rect 85580 37952 85632 38004
rect 86500 37952 86552 38004
rect 88340 37952 88392 38004
rect 88892 37952 88944 38004
rect 91744 37952 91796 38004
rect 105544 38020 105596 38072
rect 130752 38020 130804 38072
rect 141424 38020 141476 38072
rect 142160 38020 142212 38072
rect 142620 38020 142672 38072
rect 154672 38020 154724 38072
rect 155132 38020 155184 38072
rect 165620 38020 165672 38072
rect 166172 38020 166224 38072
rect 199476 38020 199528 38072
rect 328736 38020 328788 38072
rect 330484 38020 330536 38072
rect 332600 38020 332652 38072
rect 335360 38020 335412 38072
rect 336280 38020 336332 38072
rect 340144 38020 340196 38072
rect 340880 38020 340932 38072
rect 341064 38020 341116 38072
rect 369124 38020 369176 38072
rect 382832 38020 382884 38072
rect 392584 38020 392636 38072
rect 395896 38020 395948 38072
rect 460940 38020 460992 38072
rect 104164 37952 104216 38004
rect 106280 37952 106332 38004
rect 115848 37952 115900 38004
rect 116584 37952 116636 38004
rect 124220 37952 124272 38004
rect 124772 37952 124824 38004
rect 128268 37952 128320 38004
rect 129004 37952 129056 38004
rect 132132 37952 132184 38004
rect 146944 37952 146996 38004
rect 148784 37952 148836 38004
rect 217324 37952 217376 38004
rect 218796 37952 218848 38004
rect 10324 37884 10376 37936
rect 121644 37884 121696 37936
rect 136272 37884 136324 37936
rect 177304 37884 177356 37936
rect 186964 37884 187016 37936
rect 75184 37816 75236 37868
rect 77852 37816 77904 37868
rect 149520 37816 149572 37868
rect 150624 37816 150676 37868
rect 204168 37816 204220 37868
rect 206928 37816 206980 37868
rect 219440 37816 219492 37868
rect 219992 37816 220044 37868
rect 222108 37816 222160 37868
rect 222660 37816 222712 37868
rect 224224 37816 224276 37868
rect 224960 37816 225012 37868
rect 242164 37816 242216 37868
rect 242900 37816 242952 37868
rect 244924 37816 244976 37868
rect 245752 37816 245804 37868
rect 248420 37816 248472 37868
rect 248880 37816 248932 37868
rect 252560 37816 252612 37868
rect 253572 37816 253624 37868
rect 261116 37816 261168 37868
rect 262864 37816 262916 37868
rect 266360 37816 266412 37868
rect 266820 37816 266872 37868
rect 284300 37816 284352 37868
rect 284760 37816 284812 37868
rect 288440 37816 288492 37868
rect 289452 37816 289504 37868
rect 294052 37816 294104 37868
rect 294972 37816 295024 37868
rect 308036 37816 308088 37868
rect 309784 37816 309836 37868
rect 320180 37816 320232 37868
rect 320732 37816 320784 37868
rect 322204 37816 322256 37868
rect 323032 37816 323084 37868
rect 325700 37816 325752 37868
rect 326160 37816 326212 37868
rect 328736 37816 328788 37868
rect 331864 37816 331916 37868
rect 348424 37816 348476 37868
rect 350540 37816 350592 37868
rect 293132 37748 293184 37800
rect 295984 37748 296036 37800
rect 356704 37952 356756 38004
rect 358912 37952 358964 38004
rect 365720 37952 365772 38004
rect 366732 37952 366784 38004
rect 385040 37952 385092 38004
rect 385500 37952 385552 38004
rect 389180 37952 389232 38004
rect 390100 37952 390152 38004
rect 397736 37952 397788 38004
rect 467840 37952 467892 38004
rect 360844 37816 360896 37868
rect 393964 37884 394016 37936
rect 399300 37884 399352 37936
rect 474740 37884 474792 37936
rect 420920 37816 420972 37868
rect 421380 37816 421432 37868
rect 131580 37612 131632 37664
rect 133788 37612 133840 37664
rect 189172 37612 189224 37664
rect 190644 37612 190696 37664
rect 279056 37612 279108 37664
rect 280804 37612 280856 37664
rect 106280 37340 106332 37392
rect 113272 37340 113324 37392
rect 110420 37272 110472 37324
rect 114008 37272 114060 37324
rect 275192 37272 275244 37324
rect 315028 37272 315080 37324
rect 318064 37272 318116 37324
rect 353944 37272 353996 37324
rect 355048 37272 355100 37324
rect 364340 36932 364392 36984
rect 223580 36864 223632 36916
rect 343548 36864 343600 36916
rect 167460 36796 167512 36848
rect 327080 36796 327132 36848
rect 154580 36728 154632 36780
rect 228548 36728 228600 36780
rect 297824 36728 297876 36780
rect 466460 36728 466512 36780
rect 156512 36660 156564 36712
rect 277400 36660 277452 36712
rect 313188 36660 313240 36712
rect 538220 36660 538272 36712
rect 4804 36592 4856 36644
rect 41420 36592 41472 36644
rect 56508 36592 56560 36644
rect 76104 36592 76156 36644
rect 92388 36592 92440 36644
rect 122840 36592 122892 36644
rect 217876 36592 217928 36644
rect 557540 36592 557592 36644
rect 17224 36524 17276 36576
rect 93952 36524 94004 36576
rect 133788 36524 133840 36576
rect 164240 36524 164292 36576
rect 186228 36524 186280 36576
rect 412640 36524 412692 36576
rect 422760 36524 422812 36576
rect 579620 36524 579672 36576
rect 402980 35844 403032 35896
rect 403348 35844 403400 35896
rect 407120 35844 407172 35896
rect 408132 35844 408184 35896
rect 222384 35572 222436 35624
rect 243360 35572 243412 35624
rect 251180 35572 251232 35624
rect 349528 35572 349580 35624
rect 204260 35504 204312 35556
rect 239404 35504 239456 35556
rect 290096 35504 290148 35556
rect 434720 35504 434772 35556
rect 167000 35436 167052 35488
rect 330392 35436 330444 35488
rect 171416 35368 171468 35420
rect 349160 35368 349212 35420
rect 419724 35368 419776 35420
rect 571340 35368 571392 35420
rect 127072 35300 127124 35352
rect 222200 35300 222252 35352
rect 261208 35300 261260 35352
rect 303620 35300 303672 35352
rect 311992 35300 312044 35352
rect 534080 35300 534132 35352
rect 201500 35232 201552 35284
rect 483020 35232 483072 35284
rect 6920 35164 6972 35216
rect 41328 35164 41380 35216
rect 68928 35164 68980 35216
rect 121552 35164 121604 35216
rect 219532 35164 219584 35216
rect 564440 35164 564492 35216
rect 307024 34212 307076 34264
rect 360384 34212 360436 34264
rect 161480 34144 161532 34196
rect 230020 34144 230072 34196
rect 259460 34144 259512 34196
rect 351000 34144 351052 34196
rect 140872 34076 140924 34128
rect 225328 34076 225380 34128
rect 278320 34076 278372 34128
rect 378232 34076 378284 34128
rect 209872 34008 209924 34060
rect 340052 34008 340104 34060
rect 163688 33940 163740 33992
rect 313280 33940 313332 33992
rect 408776 33940 408828 33992
rect 521660 33940 521712 33992
rect 196072 33872 196124 33924
rect 458180 33872 458232 33924
rect 224132 33804 224184 33856
rect 489920 33804 489972 33856
rect 11060 33736 11112 33788
rect 42892 33736 42944 33788
rect 55220 33736 55272 33788
rect 75920 33736 75972 33788
rect 220820 33736 220872 33788
rect 572720 33736 572772 33788
rect 3148 33056 3200 33108
rect 38108 33056 38160 33108
rect 428648 33056 428700 33108
rect 579896 33056 579948 33108
rect 291844 32784 291896 32836
rect 357532 32784 357584 32836
rect 150624 32716 150676 32768
rect 245660 32716 245712 32768
rect 275928 32716 275980 32768
rect 367192 32716 367244 32768
rect 234620 32648 234672 32700
rect 345020 32648 345072 32700
rect 160192 32580 160244 32632
rect 295340 32580 295392 32632
rect 295984 32580 296036 32632
rect 445760 32580 445812 32632
rect 181628 32512 181680 32564
rect 394792 32512 394844 32564
rect 197452 32444 197504 32496
rect 465172 32444 465224 32496
rect 35900 32376 35952 32428
rect 47400 32376 47452 32428
rect 49884 32376 49936 32428
rect 100852 32376 100904 32428
rect 216772 32376 216824 32428
rect 554780 32376 554832 32428
rect 143632 31424 143684 31476
rect 226340 31424 226392 31476
rect 273260 31424 273312 31476
rect 353852 31424 353904 31476
rect 216680 31356 216732 31408
rect 340972 31356 341024 31408
rect 133880 31288 133932 31340
rect 223856 31288 223908 31340
rect 291752 31288 291804 31340
rect 441620 31288 441672 31340
rect 172704 31220 172756 31272
rect 345020 31220 345072 31272
rect 418252 31220 418304 31272
rect 564532 31220 564584 31272
rect 20720 31152 20772 31204
rect 44272 31152 44324 31204
rect 76012 31152 76064 31204
rect 199568 31152 199620 31204
rect 476120 31152 476172 31204
rect 44272 31016 44324 31068
rect 74632 31016 74684 31068
rect 206928 31084 206980 31136
rect 494060 31084 494112 31136
rect 222660 31016 222712 31068
rect 575480 31016 575532 31068
rect 76012 30948 76064 31000
rect 276112 29996 276164 30048
rect 371424 29996 371476 30048
rect 158720 29928 158772 29980
rect 229100 29928 229152 29980
rect 244372 29928 244424 29980
rect 347872 29928 347924 29980
rect 205640 29860 205692 29912
rect 339500 29860 339552 29912
rect 405740 29860 405792 29912
rect 506480 29860 506532 29912
rect 168380 29792 168432 29844
rect 334164 29792 334216 29844
rect 417424 29792 417476 29844
rect 560300 29792 560352 29844
rect 154764 29724 154816 29776
rect 270500 29724 270552 29776
rect 309600 29724 309652 29776
rect 523040 29724 523092 29776
rect 33140 29656 33192 29708
rect 46940 29656 46992 29708
rect 190644 29656 190696 29708
rect 426440 29656 426492 29708
rect 15844 29588 15896 29640
rect 92664 29588 92716 29640
rect 205088 29588 205140 29640
rect 500960 29588 501012 29640
rect 262772 28704 262824 28756
rect 310520 28704 310572 28756
rect 262220 28636 262272 28688
rect 352012 28636 352064 28688
rect 279240 28568 279292 28620
rect 385224 28568 385276 28620
rect 165712 28500 165764 28552
rect 320364 28500 320416 28552
rect 176752 28432 176804 28484
rect 333060 28432 333112 28484
rect 404452 28432 404504 28484
rect 499580 28432 499632 28484
rect 151820 28364 151872 28416
rect 259644 28364 259696 28416
rect 309784 28364 309836 28416
rect 513380 28364 513432 28416
rect 183928 28296 183980 28348
rect 405740 28296 405792 28348
rect 415768 28296 415820 28348
rect 553400 28296 553452 28348
rect 2780 28228 2832 28280
rect 66904 28228 66956 28280
rect 209044 28228 209096 28280
rect 507860 28228 507912 28280
rect 293960 27344 294012 27396
rect 356704 27344 356756 27396
rect 273720 27276 273772 27328
rect 360200 27276 360252 27328
rect 294144 27208 294196 27260
rect 452660 27208 452712 27260
rect 167552 27140 167604 27192
rect 331220 27140 331272 27192
rect 140044 27072 140096 27124
rect 323768 27072 323820 27124
rect 412824 27072 412876 27124
rect 539600 27072 539652 27124
rect 67824 27004 67876 27056
rect 104072 27004 104124 27056
rect 153568 27004 153620 27056
rect 267832 27004 267884 27056
rect 309140 27004 309192 27056
rect 520280 27004 520332 27056
rect 187056 26936 187108 26988
rect 419540 26936 419592 26988
rect 14464 26868 14516 26920
rect 67640 26868 67692 26920
rect 207388 26868 207440 26920
rect 512000 26868 512052 26920
rect 151820 25916 151872 25968
rect 227812 25916 227864 25968
rect 248604 25916 248656 25968
rect 330576 25916 330628 25968
rect 201500 25848 201552 25900
rect 338212 25848 338264 25900
rect 143724 25780 143776 25832
rect 220820 25780 220872 25832
rect 294052 25780 294104 25832
rect 456892 25780 456944 25832
rect 218704 25712 218756 25764
rect 390652 25712 390704 25764
rect 421012 25712 421064 25764
rect 574100 25712 574152 25764
rect 158812 25644 158864 25696
rect 292580 25644 292632 25696
rect 314660 25644 314712 25696
rect 547880 25644 547932 25696
rect 193220 25576 193272 25628
rect 451280 25576 451332 25628
rect 17960 25508 18012 25560
rect 69020 25508 69072 25560
rect 77300 25508 77352 25560
rect 106372 25508 106424 25560
rect 214012 25508 214064 25560
rect 543740 25508 543792 25560
rect 149060 24488 149112 24540
rect 249984 24488 250036 24540
rect 276020 24488 276072 24540
rect 353944 24488 353996 24540
rect 241612 24420 241664 24472
rect 346492 24420 346544 24472
rect 184940 24352 184992 24404
rect 333980 24352 334032 24404
rect 182180 24284 182232 24336
rect 398932 24284 398984 24336
rect 412732 24284 412784 24336
rect 542360 24284 542412 24336
rect 170404 24216 170456 24268
rect 309140 24216 309192 24268
rect 318800 24216 318852 24268
rect 565820 24216 565872 24268
rect 70584 24148 70636 24200
rect 104900 24148 104952 24200
rect 197360 24148 197412 24200
rect 469220 24148 469272 24200
rect 22100 24080 22152 24132
rect 70492 24080 70544 24132
rect 209964 24080 210016 24132
rect 523132 24080 523184 24132
rect 263784 23196 263836 23248
rect 314660 23196 314712 23248
rect 266544 23128 266596 23180
rect 351920 23128 351972 23180
rect 288532 23060 288584 23112
rect 427820 23060 427872 23112
rect 194692 22992 194744 23044
rect 336740 22992 336792 23044
rect 165620 22924 165672 22976
rect 324320 22924 324372 22976
rect 407212 22924 407264 22976
rect 514760 22924 514812 22976
rect 151912 22856 151964 22908
rect 263692 22856 263744 22908
rect 307760 22856 307812 22908
rect 516140 22856 516192 22908
rect 34520 22788 34572 22840
rect 71872 22788 71924 22840
rect 188344 22788 188396 22840
rect 408500 22788 408552 22840
rect 418160 22788 418212 22840
rect 567200 22788 567252 22840
rect 63592 22720 63644 22772
rect 103520 22720 103572 22772
rect 205732 22720 205784 22772
rect 505100 22720 505152 22772
rect 294604 21836 294656 21888
rect 357440 21836 357492 21888
rect 280804 21768 280856 21820
rect 382372 21768 382424 21820
rect 219532 21700 219584 21752
rect 342260 21700 342312 21752
rect 262312 21632 262364 21684
rect 307760 21632 307812 21684
rect 312544 21632 312596 21684
rect 463700 21632 463752 21684
rect 164332 21564 164384 21616
rect 316224 21564 316276 21616
rect 150532 21496 150584 21548
rect 256884 21496 256936 21548
rect 306380 21496 306432 21548
rect 509240 21496 509292 21548
rect 27620 21428 27672 21480
rect 70400 21428 70452 21480
rect 183560 21428 183612 21480
rect 401692 21428 401744 21480
rect 409972 21428 410024 21480
rect 528560 21428 528612 21480
rect 56784 21360 56836 21412
rect 101404 21360 101456 21412
rect 129740 21360 129792 21412
rect 157340 21360 157392 21412
rect 204352 21360 204404 21412
rect 498200 21360 498252 21412
rect 3424 20612 3476 20664
rect 38016 20612 38068 20664
rect 428556 20612 428608 20664
rect 579896 20612 579948 20664
rect 267924 20340 267976 20392
rect 332600 20340 332652 20392
rect 307116 20272 307168 20324
rect 374184 20272 374236 20324
rect 237564 20204 237616 20256
rect 346400 20204 346452 20256
rect 200764 20136 200816 20188
rect 338212 20136 338264 20188
rect 409880 20136 409932 20188
rect 524420 20136 524472 20188
rect 157524 20068 157576 20120
rect 284484 20068 284536 20120
rect 288440 20068 288492 20120
rect 432052 20068 432104 20120
rect 52644 20000 52696 20052
rect 76012 20000 76064 20052
rect 189080 20000 189132 20052
rect 430580 20000 430632 20052
rect 74632 19932 74684 19984
rect 104164 19932 104216 19984
rect 139492 19932 139544 19984
rect 207020 19932 207072 19984
rect 215300 19932 215352 19984
rect 550640 19932 550692 19984
rect 255504 18980 255556 19032
rect 348424 18980 348476 19032
rect 139400 18912 139452 18964
rect 202880 18912 202932 18964
rect 280252 18912 280304 18964
rect 389364 18912 389416 18964
rect 174084 18844 174136 18896
rect 330484 18844 330536 18896
rect 172612 18776 172664 18828
rect 351920 18776 351972 18828
rect 407120 18776 407172 18828
rect 517520 18776 517572 18828
rect 157432 18708 157484 18760
rect 288440 18708 288492 18760
rect 310612 18708 310664 18760
rect 527180 18708 527232 18760
rect 48320 18640 48372 18692
rect 74540 18640 74592 18692
rect 195244 18640 195296 18692
rect 448520 18640 448572 18692
rect 60924 18572 60976 18624
rect 102232 18572 102284 18624
rect 201592 18572 201644 18624
rect 487160 18572 487212 18624
rect 269304 17620 269356 17672
rect 353300 17620 353352 17672
rect 212724 17552 212776 17604
rect 340144 17552 340196 17604
rect 136824 17484 136876 17536
rect 224224 17484 224276 17536
rect 291200 17484 291252 17536
rect 438860 17484 438912 17536
rect 169760 17416 169812 17468
rect 340972 17416 341024 17468
rect 416780 17416 416832 17468
rect 556160 17416 556212 17468
rect 195980 17348 196032 17400
rect 462320 17348 462372 17400
rect 66260 17280 66312 17332
rect 78772 17280 78824 17332
rect 200120 17280 200172 17332
rect 480260 17280 480312 17332
rect 8300 17212 8352 17264
rect 67732 17212 67784 17264
rect 88432 17212 88484 17264
rect 104900 17212 104952 17264
rect 134064 17212 134116 17264
rect 182180 17212 182232 17264
rect 219440 17212 219492 17264
rect 568580 17212 568632 17264
rect 298284 16396 298336 16448
rect 358912 16396 358964 16448
rect 227536 16328 227588 16380
rect 343732 16328 343784 16380
rect 198740 16260 198792 16312
rect 338120 16260 338172 16312
rect 331864 16192 331916 16244
rect 473452 16192 473504 16244
rect 192024 16124 192076 16176
rect 335360 16124 335412 16176
rect 188528 16056 188580 16108
rect 335452 16056 335504 16108
rect 292672 15988 292724 16040
rect 448612 15988 448664 16040
rect 81624 15920 81676 15972
rect 107752 15920 107804 15972
rect 133972 15920 134024 15972
rect 178592 15920 178644 15972
rect 180984 15920 181036 15972
rect 334072 15920 334124 15972
rect 342904 15920 342956 15972
rect 547972 15920 548024 15972
rect 59360 15852 59412 15904
rect 93952 15852 94004 15904
rect 147864 15852 147916 15904
rect 226432 15852 226484 15904
rect 318064 15852 318116 15904
rect 545488 15852 545540 15904
rect 262864 14968 262916 15020
rect 300768 14968 300820 15020
rect 280712 14900 280764 14952
rect 356152 14900 356204 14952
rect 231032 14832 231084 14884
rect 345112 14832 345164 14884
rect 170312 14764 170364 14816
rect 331312 14764 331364 14816
rect 218060 14696 218112 14748
rect 242164 14696 242216 14748
rect 295432 14696 295484 14748
rect 459928 14696 459980 14748
rect 211712 14628 211764 14680
rect 240232 14628 240284 14680
rect 298192 14628 298244 14680
rect 470600 14628 470652 14680
rect 193220 14560 193272 14612
rect 237472 14560 237524 14612
rect 298100 14560 298152 14612
rect 474096 14560 474148 14612
rect 30840 14492 30892 14544
rect 71780 14492 71832 14544
rect 129004 14492 129056 14544
rect 150624 14492 150676 14544
rect 155960 14492 156012 14544
rect 281724 14492 281776 14544
rect 299572 14492 299624 14544
rect 478144 14492 478196 14544
rect 64972 14424 65024 14476
rect 114744 14424 114796 14476
rect 129096 14424 129148 14476
rect 321560 14424 321612 14476
rect 414020 14424 414072 14476
rect 546500 14424 546552 14476
rect 280160 13676 280212 13728
rect 392492 13676 392544 13728
rect 281540 13608 281592 13660
rect 396172 13608 396224 13660
rect 281632 13540 281684 13592
rect 400128 13540 400180 13592
rect 217324 13472 217376 13524
rect 242900 13472 242952 13524
rect 282920 13472 282972 13524
rect 403624 13472 403676 13524
rect 404360 13472 404412 13524
rect 503720 13472 503772 13524
rect 215300 13404 215352 13456
rect 241520 13404 241572 13456
rect 284392 13404 284444 13456
rect 407120 13404 407172 13456
rect 132592 13336 132644 13388
rect 175464 13336 175516 13388
rect 201592 13336 201644 13388
rect 238760 13336 238812 13388
rect 284300 13336 284352 13388
rect 410800 13336 410852 13388
rect 411260 13336 411312 13388
rect 536104 13336 536156 13388
rect 166080 13268 166132 13320
rect 230480 13268 230532 13320
rect 285772 13268 285824 13320
rect 417424 13268 417476 13320
rect 154672 13200 154724 13252
rect 274824 13200 274876 13252
rect 287152 13200 287204 13252
rect 421012 13200 421064 13252
rect 63500 13132 63552 13184
rect 111616 13132 111668 13184
rect 163688 13132 163740 13184
rect 286324 13132 286376 13184
rect 287060 13132 287112 13184
rect 424968 13132 425020 13184
rect 30104 13064 30156 13116
rect 45560 13064 45612 13116
rect 53288 13064 53340 13116
rect 100760 13064 100812 13116
rect 138848 13064 138900 13116
rect 282184 13064 282236 13116
rect 285680 13064 285732 13116
rect 414296 13064 414348 13116
rect 414664 13064 414716 13116
rect 576952 13064 577004 13116
rect 249892 12316 249944 12368
rect 254216 12316 254268 12368
rect 197912 12248 197964 12300
rect 237380 12248 237432 12300
rect 266452 12248 266504 12300
rect 324412 12248 324464 12300
rect 190644 12180 190696 12232
rect 236000 12180 236052 12232
rect 266360 12180 266412 12232
rect 328736 12180 328788 12232
rect 186872 12112 186924 12164
rect 234712 12112 234764 12164
rect 267740 12112 267792 12164
rect 336280 12112 336332 12164
rect 183744 12044 183796 12096
rect 234804 12044 234856 12096
rect 269212 12044 269264 12096
rect 339500 12044 339552 12096
rect 180248 11976 180300 12028
rect 233332 11976 233384 12028
rect 269120 11976 269172 12028
rect 342904 11976 342956 12028
rect 393964 11976 394016 12028
rect 415492 11976 415544 12028
rect 176844 11908 176896 11960
rect 233240 11908 233292 11960
rect 270592 11908 270644 11960
rect 346952 11908 347004 11960
rect 383660 11908 383712 11960
rect 407212 11908 407264 11960
rect 172704 11840 172756 11892
rect 231952 11840 232004 11892
rect 249800 11840 249852 11892
rect 251456 11840 251508 11892
rect 271880 11840 271932 11892
rect 353576 11840 353628 11892
rect 405832 11840 405884 11892
rect 511264 11840 511316 11892
rect 37832 11772 37884 11824
rect 71044 11772 71096 11824
rect 85672 11772 85724 11824
rect 107660 11772 107712 11824
rect 168380 11772 168432 11824
rect 231860 11772 231912 11824
rect 236552 11772 236604 11824
rect 245752 11772 245804 11824
rect 270684 11772 270736 11824
rect 349252 11772 349304 11824
rect 349804 11772 349856 11824
rect 531320 11772 531372 11824
rect 60832 11704 60884 11756
rect 100760 11704 100812 11756
rect 105544 11704 105596 11756
rect 119896 11704 119948 11756
rect 130568 11704 130620 11756
rect 222292 11704 222344 11756
rect 233424 11704 233476 11756
rect 244924 11704 244976 11756
rect 273352 11704 273404 11756
rect 357532 11704 357584 11756
rect 360844 11704 360896 11756
rect 562048 11704 562100 11756
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 423680 11568 423732 11620
rect 240232 11364 240284 11416
rect 247040 11364 247092 11416
rect 423772 11364 423824 11416
rect 187700 10616 187752 10668
rect 423864 10616 423916 10668
rect 425704 10616 425756 10668
rect 532056 10616 532108 10668
rect 190552 10548 190604 10600
rect 433984 10548 434036 10600
rect 436744 10548 436796 10600
rect 550272 10548 550324 10600
rect 190460 10480 190512 10532
rect 437480 10480 437532 10532
rect 191932 10412 191984 10464
rect 440332 10412 440384 10464
rect 41880 10344 41932 10396
rect 72424 10344 72476 10396
rect 89720 10344 89772 10396
rect 112352 10344 112404 10396
rect 191840 10344 191892 10396
rect 445024 10344 445076 10396
rect 17040 10276 17092 10328
rect 42800 10276 42852 10328
rect 60740 10276 60792 10328
rect 97448 10276 97500 10328
rect 132500 10276 132552 10328
rect 171968 10276 172020 10328
rect 177304 10276 177356 10328
rect 186136 10276 186188 10328
rect 194600 10276 194652 10328
rect 455696 10276 455748 10328
rect 172520 9528 172572 9580
rect 356336 9528 356388 9580
rect 173992 9460 174044 9512
rect 359924 9460 359976 9512
rect 173900 9392 173952 9444
rect 363512 9392 363564 9444
rect 175280 9324 175332 9376
rect 367008 9324 367060 9376
rect 175372 9256 175424 9308
rect 370596 9256 370648 9308
rect 382280 9256 382332 9308
rect 404820 9256 404872 9308
rect 176660 9188 176712 9240
rect 374092 9188 374144 9240
rect 380992 9188 381044 9240
rect 397736 9188 397788 9240
rect 400220 9188 400272 9240
rect 482836 9188 482888 9240
rect 178040 9120 178092 9172
rect 377680 9120 377732 9172
rect 400312 9120 400364 9172
rect 486424 9120 486476 9172
rect 85764 9052 85816 9104
rect 95148 9052 95200 9104
rect 178132 9052 178184 9104
rect 381176 9052 381228 9104
rect 401600 9052 401652 9104
rect 489920 9052 489972 9104
rect 53932 8984 53984 9036
rect 69112 8984 69164 9036
rect 70308 8984 70360 9036
rect 80152 8984 80204 9036
rect 87052 8984 87104 9036
rect 102232 8984 102284 9036
rect 146944 8984 146996 9036
rect 168472 8984 168524 9036
rect 179420 8984 179472 9036
rect 384764 8984 384816 9036
rect 403072 8984 403124 9036
rect 493508 8984 493560 9036
rect 3976 8916 4028 8968
rect 40132 8916 40184 8968
rect 63224 8916 63276 8968
rect 78680 8916 78732 8968
rect 93124 8916 93176 8968
rect 116400 8916 116452 8968
rect 128360 8916 128412 8968
rect 154212 8916 154264 8968
rect 179512 8916 179564 8968
rect 388260 8916 388312 8968
rect 392584 8916 392636 8968
rect 401324 8916 401376 8968
rect 402980 8916 403032 8968
rect 497096 8916 497148 8968
rect 80888 8712 80940 8764
rect 82912 8712 82964 8764
rect 284300 8168 284352 8220
rect 324964 8168 325016 8220
rect 263600 8100 263652 8152
rect 318524 8100 318576 8152
rect 131764 8032 131816 8084
rect 322204 8032 322256 8084
rect 313372 7964 313424 8016
rect 541992 7964 542044 8016
rect 316040 7896 316092 7948
rect 552664 7896 552716 7948
rect 316132 7828 316184 7880
rect 556160 7828 556212 7880
rect 208584 7760 208636 7812
rect 240140 7760 240192 7812
rect 259552 7760 259604 7812
rect 297272 7760 297324 7812
rect 317420 7760 317472 7812
rect 559748 7760 559800 7812
rect 85580 7692 85632 7744
rect 98644 7692 98696 7744
rect 160100 7692 160152 7744
rect 299664 7692 299716 7744
rect 317512 7692 317564 7744
rect 563244 7692 563296 7744
rect 53840 7624 53892 7676
rect 65524 7624 65576 7676
rect 69664 7624 69716 7676
rect 90364 7624 90416 7676
rect 161664 7624 161716 7676
rect 303160 7624 303212 7676
rect 320272 7624 320324 7676
rect 570328 7624 570380 7676
rect 26516 7556 26568 7608
rect 44180 7556 44232 7608
rect 59636 7556 59688 7608
rect 75184 7556 75236 7608
rect 88340 7556 88392 7608
rect 109316 7556 109368 7608
rect 141424 7556 141476 7608
rect 161296 7556 161348 7608
rect 161572 7556 161624 7608
rect 306748 7556 306800 7608
rect 320180 7556 320232 7608
rect 573916 7556 573968 7608
rect 218060 7488 218112 7540
rect 219256 7488 219308 7540
rect 77392 7216 77444 7268
rect 81440 7216 81492 7268
rect 3424 6808 3476 6860
rect 37924 6808 37976 6860
rect 252652 6808 252704 6860
rect 265348 6808 265400 6860
rect 428556 6808 428608 6860
rect 580172 6808 580224 6860
rect 264980 6672 265032 6724
rect 322112 6672 322164 6724
rect 251364 6604 251416 6656
rect 261760 6604 261812 6656
rect 299480 6604 299532 6656
rect 481732 6604 481784 6656
rect 252560 6536 252612 6588
rect 268844 6536 268896 6588
rect 300860 6536 300912 6588
rect 485228 6536 485280 6588
rect 143540 6468 143592 6520
rect 225144 6468 225196 6520
rect 253940 6468 253992 6520
rect 272432 6468 272484 6520
rect 302240 6468 302292 6520
rect 488816 6468 488868 6520
rect 144920 6400 144972 6452
rect 228732 6400 228784 6452
rect 229836 6400 229888 6452
rect 244464 6400 244516 6452
rect 255412 6400 255464 6452
rect 276020 6400 276072 6452
rect 302332 6400 302384 6452
rect 492312 6400 492364 6452
rect 145012 6332 145064 6384
rect 232228 6332 232280 6384
rect 255320 6332 255372 6384
rect 279516 6332 279568 6384
rect 303804 6332 303856 6384
rect 495900 6332 495952 6384
rect 146300 6264 146352 6316
rect 235816 6264 235868 6316
rect 256700 6264 256752 6316
rect 283104 6264 283156 6316
rect 303712 6264 303764 6316
rect 499396 6264 499448 6316
rect 58624 6196 58676 6248
rect 72608 6196 72660 6248
rect 73804 6196 73856 6248
rect 80060 6196 80112 6248
rect 147680 6196 147732 6248
rect 239312 6196 239364 6248
rect 256792 6196 256844 6248
rect 286600 6196 286652 6248
rect 305000 6196 305052 6248
rect 502984 6196 503036 6248
rect 52552 6128 52604 6180
rect 58440 6128 58492 6180
rect 64880 6128 64932 6180
rect 118792 6128 118844 6180
rect 150440 6128 150492 6180
rect 253480 6128 253532 6180
rect 258172 6128 258224 6180
rect 293684 6128 293736 6180
rect 305092 6128 305144 6180
rect 506480 6128 506532 6180
rect 244096 5584 244148 5636
rect 248512 5584 248564 5636
rect 44272 5516 44324 5568
rect 46204 5516 46256 5568
rect 84200 5516 84252 5568
rect 91560 5516 91612 5568
rect 247592 5516 247644 5568
rect 248420 5516 248472 5568
rect 142252 5312 142304 5364
rect 214472 5312 214524 5364
rect 142160 5244 142212 5296
rect 218152 5244 218204 5296
rect 258080 5244 258132 5296
rect 290188 5244 290240 5296
rect 208492 5176 208544 5228
rect 515956 5176 516008 5228
rect 208400 5108 208452 5160
rect 519544 5108 519596 5160
rect 56692 5040 56744 5092
rect 79692 5040 79744 5092
rect 136732 5040 136784 5092
rect 189724 5040 189776 5092
rect 209780 5040 209832 5092
rect 526628 5040 526680 5092
rect 56600 4972 56652 5024
rect 83280 4972 83332 5024
rect 136640 4972 136692 5024
rect 193312 4972 193364 5024
rect 211160 4972 211212 5024
rect 530124 4972 530176 5024
rect 57980 4904 58032 4956
rect 86868 4904 86920 4956
rect 138020 4904 138072 4956
rect 196808 4904 196860 4956
rect 212632 4904 212684 4956
rect 533712 4904 533764 4956
rect 62212 4836 62264 4888
rect 104532 4836 104584 4888
rect 138112 4836 138164 4888
rect 200304 4836 200356 4888
rect 212540 4836 212592 4888
rect 537208 4836 537260 4888
rect 572 4768 624 4820
rect 39304 4768 39356 4820
rect 52460 4768 52512 4820
rect 62028 4768 62080 4820
rect 62120 4768 62172 4820
rect 108120 4768 108172 4820
rect 140780 4768 140832 4820
rect 210976 4768 211028 4820
rect 213920 4700 213972 4752
rect 540796 4768 540848 4820
rect 40684 4564 40736 4616
rect 47584 4564 47636 4616
rect 251272 4496 251324 4548
rect 258264 4496 258316 4548
rect 82820 4292 82872 4344
rect 84476 4292 84528 4344
rect 49700 4224 49752 4276
rect 51356 4224 51408 4276
rect 47860 4156 47912 4208
rect 49792 4156 49844 4208
rect 51080 4156 51132 4208
rect 54944 4156 54996 4208
rect 14740 4088 14792 4140
rect 17224 4088 17276 4140
rect 43076 4088 43128 4140
rect 98000 4088 98052 4140
rect 323308 4088 323360 4140
rect 364524 4088 364576 4140
rect 389180 4088 389232 4140
rect 436744 4088 436796 4140
rect 39580 4020 39632 4072
rect 98092 4020 98144 4072
rect 319720 4020 319772 4072
rect 364432 4020 364484 4072
rect 390560 4020 390612 4072
rect 440240 4020 440292 4072
rect 35992 3952 36044 4004
rect 96712 3952 96764 4004
rect 316224 3952 316276 4004
rect 362960 3952 363012 4004
rect 391940 3952 391992 4004
rect 443828 3952 443880 4004
rect 32404 3884 32456 3936
rect 96620 3884 96672 3936
rect 121644 3884 121696 3936
rect 125876 3884 125928 3936
rect 312636 3884 312688 3936
rect 363052 3884 363104 3936
rect 385040 3884 385092 3936
rect 392032 3884 392084 3936
rect 393320 3884 393372 3936
rect 450912 3884 450964 3936
rect 28908 3816 28960 3868
rect 95332 3816 95384 3868
rect 103336 3816 103388 3868
rect 111892 3816 111944 3868
rect 24216 3748 24268 3800
rect 95240 3748 95292 3800
rect 99840 3748 99892 3800
rect 111800 3748 111852 3800
rect 19432 3680 19484 3732
rect 94044 3680 94096 3732
rect 96252 3680 96304 3732
rect 110604 3680 110656 3732
rect 25320 3612 25372 3664
rect 120172 3816 120224 3868
rect 168380 3816 168432 3868
rect 169576 3816 169628 3868
rect 176752 3816 176804 3868
rect 177856 3816 177908 3868
rect 251180 3816 251232 3868
rect 252376 3816 252428 3868
rect 291384 3816 291436 3868
rect 294604 3816 294656 3868
rect 309048 3816 309100 3868
rect 361672 3816 361724 3868
rect 362316 3816 362368 3868
rect 374000 3816 374052 3868
rect 379520 3816 379572 3868
rect 387156 3816 387208 3868
rect 394700 3816 394752 3868
rect 458088 3816 458140 3868
rect 160100 3748 160152 3800
rect 328552 3748 328604 3800
rect 348056 3748 348108 3800
rect 369952 3748 370004 3800
rect 379612 3748 379664 3800
rect 390560 3748 390612 3800
rect 396080 3748 396132 3800
rect 465172 3748 465224 3800
rect 124312 3680 124364 3732
rect 132960 3680 133012 3732
rect 135260 3680 135312 3732
rect 140044 3680 140096 3732
rect 156604 3680 156656 3732
rect 328460 3680 328512 3732
rect 344560 3680 344612 3732
rect 369860 3680 369912 3732
rect 372896 3680 372948 3732
rect 375564 3680 375616 3732
rect 380900 3680 380952 3732
rect 394240 3680 394292 3732
rect 397460 3680 397512 3732
rect 472256 3680 472308 3732
rect 9956 3544 10008 3596
rect 15844 3544 15896 3596
rect 20628 3544 20680 3596
rect 118976 3612 119028 3664
rect 124220 3612 124272 3664
rect 136456 3612 136508 3664
rect 153016 3612 153068 3664
rect 327172 3612 327224 3664
rect 337476 3612 337528 3664
rect 368572 3612 368624 3664
rect 385132 3612 385184 3664
rect 407028 3612 407080 3664
rect 407212 3612 407264 3664
rect 408408 3612 408460 3664
rect 2872 3476 2924 3528
rect 4804 3476 4856 3528
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 15936 3476 15988 3528
rect 118700 3544 118752 3596
rect 126980 3544 127032 3596
rect 147128 3544 147180 3596
rect 149520 3544 149572 3596
rect 327264 3544 327316 3596
rect 333888 3544 333940 3596
rect 367100 3544 367152 3596
rect 386420 3544 386472 3596
rect 116584 3476 116636 3528
rect 117596 3476 117648 3528
rect 128176 3476 128228 3528
rect 129096 3476 129148 3528
rect 6460 3408 6512 3460
rect 10324 3408 10376 3460
rect 11152 3408 11204 3460
rect 117320 3408 117372 3460
rect 125600 3408 125652 3460
rect 143540 3476 143592 3528
rect 145932 3476 145984 3528
rect 325700 3476 325752 3528
rect 330392 3476 330444 3528
rect 365720 3476 365772 3528
rect 390652 3476 390704 3528
rect 391848 3476 391900 3528
rect 392032 3544 392084 3596
rect 415400 3612 415452 3664
rect 423588 3612 423640 3664
rect 582196 3612 582248 3664
rect 418988 3544 419040 3596
rect 420920 3544 420972 3596
rect 578608 3544 578660 3596
rect 415492 3476 415544 3528
rect 416688 3476 416740 3528
rect 422392 3476 422444 3528
rect 581000 3476 581052 3528
rect 46664 3340 46716 3392
rect 99380 3340 99432 3392
rect 125692 3340 125744 3392
rect 140044 3408 140096 3460
rect 142436 3408 142488 3460
rect 325792 3408 325844 3460
rect 326804 3408 326856 3460
rect 193220 3340 193272 3392
rect 194416 3340 194468 3392
rect 287796 3340 287848 3392
rect 291844 3340 291896 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 351644 3340 351696 3392
rect 365812 3408 365864 3460
rect 374184 3408 374236 3460
rect 386512 3408 386564 3460
rect 422576 3408 422628 3460
rect 423680 3408 423732 3460
rect 583392 3408 583444 3460
rect 89168 3272 89220 3324
rect 109040 3272 109092 3324
rect 116032 3272 116084 3324
rect 124680 3272 124732 3324
rect 355232 3272 355284 3324
rect 365904 3340 365956 3392
rect 389272 3340 389324 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 523040 3340 523092 3392
rect 523868 3340 523920 3392
rect 547880 3340 547932 3392
rect 548708 3340 548760 3392
rect 564440 3340 564492 3392
rect 565268 3340 565320 3392
rect 92756 3204 92808 3256
rect 109132 3204 109184 3256
rect 122932 3204 122984 3256
rect 129372 3204 129424 3256
rect 371240 3272 371292 3324
rect 376944 3272 376996 3324
rect 379980 3272 380032 3324
rect 387892 3272 387944 3324
rect 429660 3272 429712 3324
rect 371332 3204 371384 3256
rect 387800 3204 387852 3256
rect 426164 3204 426216 3256
rect 369400 3136 369452 3188
rect 375472 3136 375524 3188
rect 407028 3136 407080 3188
rect 411904 3136 411956 3188
rect 115940 3068 115992 3120
rect 121092 3068 121144 3120
rect 358728 3068 358780 3120
rect 372620 3068 372672 3120
rect 1676 3000 1728 3052
rect 3976 3000 4028 3052
rect 378140 2932 378192 2984
rect 383568 2932 383620 2984
rect 301964 2864 302016 2916
rect 307024 2864 307076 2916
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 683806 3464 697303
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3424 683800 3476 683806
rect 3424 683742 3476 683748
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2870 645144 2926 645153
rect 2870 645079 2926 645088
rect 2884 644502 2912 645079
rect 2872 644496 2924 644502
rect 2872 644438 2924 644444
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3330 593056 3386 593065
rect 3330 592991 3386 593000
rect 3344 592074 3372 592991
rect 3332 592068 3384 592074
rect 3332 592010 3384 592016
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553586 3188 553823
rect 3148 553580 3200 553586
rect 3148 553522 3200 553528
rect 3054 540832 3110 540841
rect 3054 540767 3110 540776
rect 3068 539646 3096 540767
rect 3056 539640 3108 539646
rect 3056 539582 3108 539588
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3436 527134 3464 671191
rect 3528 671022 3556 684247
rect 3516 671016 3568 671022
rect 3516 670958 3568 670964
rect 4804 671016 4856 671022
rect 4804 670958 4856 670964
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3424 527128 3476 527134
rect 3424 527070 3476 527076
rect 3422 514856 3478 514865
rect 3422 514791 3478 514800
rect 3146 488744 3202 488753
rect 3146 488679 3202 488688
rect 3160 488578 3188 488679
rect 3148 488572 3200 488578
rect 3148 488514 3200 488520
rect 3330 436656 3386 436665
rect 3330 436591 3386 436600
rect 3344 436150 3372 436591
rect 3332 436144 3384 436150
rect 3332 436086 3384 436092
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 422346 3372 423535
rect 3332 422340 3384 422346
rect 3332 422282 3384 422288
rect 3436 412622 3464 514791
rect 3528 488510 3556 619103
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 488504 3568 488510
rect 3516 488446 3568 488452
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3528 474774 3556 475623
rect 3516 474768 3568 474774
rect 3516 474710 3568 474716
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3424 412616 3476 412622
rect 3424 412558 3476 412564
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3330 384432 3386 384441
rect 3330 384367 3386 384376
rect 3344 383722 3372 384367
rect 3332 383716 3384 383722
rect 3332 383658 3384 383664
rect 3146 371376 3202 371385
rect 3146 371311 3148 371320
rect 3200 371311 3202 371320
rect 3148 371282 3200 371288
rect 3436 336734 3464 410479
rect 3528 373998 3556 462567
rect 3620 449886 3648 566879
rect 4816 536790 4844 670958
rect 6932 562358 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 11704 683800 11756 683806
rect 11704 683742 11756 683748
rect 10324 644496 10376 644502
rect 10324 644438 10376 644444
rect 6920 562352 6972 562358
rect 6920 562294 6972 562300
rect 6184 553580 6236 553586
rect 6184 553522 6236 553528
rect 4804 536784 4856 536790
rect 4804 536726 4856 536732
rect 3698 501800 3754 501809
rect 3698 501735 3754 501744
rect 3608 449880 3660 449886
rect 3608 449822 3660 449828
rect 3712 402966 3740 501735
rect 3790 449576 3846 449585
rect 3790 449511 3846 449520
rect 3700 402960 3752 402966
rect 3700 402902 3752 402908
rect 3606 397488 3662 397497
rect 3606 397423 3662 397432
rect 3516 373992 3568 373998
rect 3516 373934 3568 373940
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3424 336728 3476 336734
rect 3424 336670 3476 336676
rect 2778 332344 2834 332353
rect 2778 332279 2834 332288
rect 2792 331634 2820 332279
rect 2780 331628 2832 331634
rect 2780 331570 2832 331576
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 269074 3464 319223
rect 3528 298110 3556 358391
rect 3620 327078 3648 397423
rect 3804 364342 3832 449511
rect 6196 441590 6224 553522
rect 10336 507822 10364 644438
rect 11716 545086 11744 683742
rect 22744 632120 22796 632126
rect 22744 632062 22796 632068
rect 14464 592068 14516 592074
rect 14464 592010 14516 592016
rect 11704 545080 11756 545086
rect 11704 545022 11756 545028
rect 10324 507816 10376 507822
rect 10324 507758 10376 507764
rect 10324 488572 10376 488578
rect 10324 488514 10376 488520
rect 6184 441584 6236 441590
rect 6184 441526 6236 441532
rect 10336 393310 10364 488514
rect 14476 469198 14504 592010
rect 22756 541686 22784 632062
rect 23492 562426 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 33784 656940 33836 656946
rect 33784 656882 33836 656888
rect 25504 579692 25556 579698
rect 25504 579634 25556 579640
rect 23480 562420 23532 562426
rect 23480 562362 23532 562368
rect 22744 541680 22796 541686
rect 22744 541622 22796 541628
rect 22744 539640 22796 539646
rect 22744 539582 22796 539588
rect 14464 469192 14516 469198
rect 14464 469134 14516 469140
rect 11704 436144 11756 436150
rect 11704 436086 11756 436092
rect 10324 393304 10376 393310
rect 10324 393246 10376 393252
rect 6184 371340 6236 371346
rect 6184 371282 6236 371288
rect 3792 364336 3844 364342
rect 3792 364278 3844 364284
rect 3698 345400 3754 345409
rect 3698 345335 3754 345344
rect 3608 327072 3660 327078
rect 3608 327014 3660 327020
rect 3606 306232 3662 306241
rect 3606 306167 3662 306176
rect 3516 298104 3568 298110
rect 3516 298046 3568 298052
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3424 269068 3476 269074
rect 3424 269010 3476 269016
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 231810 3464 267135
rect 3528 249762 3556 293111
rect 3620 259418 3648 306167
rect 3712 288386 3740 345335
rect 4804 331628 4856 331634
rect 4804 331570 4856 331576
rect 3700 288380 3752 288386
rect 3700 288322 3752 288328
rect 3698 280120 3754 280129
rect 3698 280055 3754 280064
rect 3608 259412 3660 259418
rect 3608 259354 3660 259360
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 3516 249756 3568 249762
rect 3516 249698 3568 249704
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3424 231804 3476 231810
rect 3424 231746 3476 231752
rect 3422 228032 3478 228041
rect 3422 227967 3478 227976
rect 3436 202842 3464 227967
rect 3528 212498 3556 241023
rect 3620 222154 3648 254079
rect 3712 240106 3740 280055
rect 4816 278730 4844 331570
rect 6196 307766 6224 371282
rect 11716 354686 11744 436086
rect 22756 431934 22784 539582
rect 25516 459542 25544 579634
rect 28264 527196 28316 527202
rect 28264 527138 28316 527144
rect 25504 459536 25556 459542
rect 25504 459478 25556 459484
rect 22744 431928 22796 431934
rect 22744 431870 22796 431876
rect 26884 422340 26936 422346
rect 26884 422282 26936 422288
rect 24124 383716 24176 383722
rect 24124 383658 24176 383664
rect 11704 354680 11756 354686
rect 11704 354622 11756 354628
rect 24136 317422 24164 383658
rect 26896 345030 26924 422282
rect 28276 422278 28304 527138
rect 33796 517478 33824 656882
rect 36544 605872 36596 605878
rect 36544 605814 36596 605820
rect 33784 517472 33836 517478
rect 33784 517414 33836 517420
rect 36556 478417 36584 605814
rect 40052 562494 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 56796 683114 56824 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 56612 683086 56824 683114
rect 40040 562488 40092 562494
rect 40040 562430 40092 562436
rect 50620 562420 50672 562426
rect 50620 562362 50672 562368
rect 40408 562352 40460 562358
rect 40408 562294 40460 562300
rect 40420 559042 40448 562294
rect 50632 559042 50660 562362
rect 56612 562358 56640 683086
rect 71792 562494 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 563038 88380 702406
rect 88340 563032 88392 563038
rect 88340 562974 88392 562980
rect 94596 563032 94648 563038
rect 94596 562974 94648 562980
rect 61660 562488 61712 562494
rect 61660 562430 61712 562436
rect 71780 562488 71832 562494
rect 71780 562430 71832 562436
rect 83648 562488 83700 562494
rect 83648 562430 83700 562436
rect 56600 562352 56652 562358
rect 56600 562294 56652 562300
rect 61672 559042 61700 562430
rect 72700 562352 72752 562358
rect 72700 562294 72752 562300
rect 72712 559042 72740 562294
rect 83660 559042 83688 562430
rect 94608 559042 94636 562974
rect 104912 559042 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 121656 699718 121684 703520
rect 137848 700330 137876 703520
rect 149060 700392 149112 700398
rect 149060 700334 149112 700340
rect 126980 700324 127032 700330
rect 126980 700266 127032 700272
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 138020 700324 138072 700330
rect 138020 700266 138072 700272
rect 115940 699712 115992 699718
rect 115940 699654 115992 699660
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 115952 559042 115980 699654
rect 126992 559042 127020 700266
rect 138032 559042 138060 700266
rect 149072 559042 149100 700334
rect 154132 700330 154160 703520
rect 170324 700398 170352 703520
rect 171140 700460 171192 700466
rect 171140 700402 171192 700408
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 160100 700324 160152 700330
rect 160100 700266 160152 700272
rect 160112 559042 160140 700266
rect 171152 559042 171180 700402
rect 182180 700392 182232 700398
rect 182180 700334 182232 700340
rect 182192 559042 182220 700334
rect 186516 700330 186544 703520
rect 202800 700466 202828 703520
rect 204260 700528 204312 700534
rect 204260 700470 204312 700476
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 186504 700324 186556 700330
rect 186504 700266 186556 700272
rect 193220 700324 193272 700330
rect 193220 700266 193272 700272
rect 193232 559042 193260 700266
rect 204272 559042 204300 700470
rect 215300 700460 215352 700466
rect 215300 700402 215352 700408
rect 215312 559042 215340 700402
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 226340 700392 226392 700398
rect 226340 700334 226392 700340
rect 226352 559042 226380 700334
rect 235184 700330 235212 703520
rect 248420 700664 248472 700670
rect 248420 700606 248472 700612
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 237380 700324 237432 700330
rect 237380 700266 237432 700272
rect 237392 559042 237420 700266
rect 248432 559042 248460 700606
rect 251468 700534 251496 703520
rect 259460 700596 259512 700602
rect 259460 700538 259512 700544
rect 251456 700528 251508 700534
rect 251456 700470 251508 700476
rect 259472 559042 259500 700538
rect 267660 700466 267688 703520
rect 270500 700528 270552 700534
rect 270500 700470 270552 700476
rect 267648 700460 267700 700466
rect 267648 700402 267700 700408
rect 270512 559042 270540 700470
rect 281540 700460 281592 700466
rect 281540 700402 281592 700408
rect 281552 559042 281580 700402
rect 283852 700398 283880 703520
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 292580 700392 292632 700398
rect 292580 700334 292632 700340
rect 292592 559042 292620 700334
rect 300136 700330 300164 703520
rect 314660 701004 314712 701010
rect 314660 700946 314712 700952
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 303620 700324 303672 700330
rect 303620 700266 303672 700272
rect 303632 559042 303660 700266
rect 314672 559042 314700 700946
rect 316328 700670 316356 703520
rect 325700 700936 325752 700942
rect 325700 700878 325752 700884
rect 316316 700664 316368 700670
rect 316316 700606 316368 700612
rect 325712 559042 325740 700878
rect 332520 700602 332548 703520
rect 336740 700868 336792 700874
rect 336740 700810 336792 700816
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 336752 559042 336780 700810
rect 347872 700800 347924 700806
rect 347872 700742 347924 700748
rect 347884 559314 347912 700742
rect 348804 700534 348832 703520
rect 358820 700732 358872 700738
rect 358820 700674 358872 700680
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 347846 559286 347912 559314
rect 40420 559014 40740 559042
rect 50632 559014 50980 559042
rect 61672 559014 61960 559042
rect 72712 559014 72960 559042
rect 83660 559014 83960 559042
rect 94608 559014 94940 559042
rect 104912 559014 105940 559042
rect 115952 559014 116940 559042
rect 126992 559014 127940 559042
rect 138032 559014 138920 559042
rect 149072 559014 149920 559042
rect 160112 559014 160920 559042
rect 171152 559014 171920 559042
rect 182192 559014 182900 559042
rect 193232 559014 193900 559042
rect 204272 559014 204920 559042
rect 215312 559014 215920 559042
rect 226352 559014 226920 559042
rect 237392 559014 237900 559042
rect 248432 559014 248900 559042
rect 259472 559014 259900 559042
rect 270512 559014 270900 559042
rect 281552 559014 281880 559042
rect 292592 559014 292880 559042
rect 303632 559014 303880 559042
rect 314672 559014 314880 559042
rect 325712 559014 325860 559042
rect 336752 559014 336860 559042
rect 347846 559028 347874 559286
rect 358832 559014 358860 700674
rect 364996 700466 365024 703520
rect 369860 700664 369912 700670
rect 369860 700606 369912 700612
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 369872 559314 369900 700606
rect 379520 700596 379572 700602
rect 379520 700538 379572 700544
rect 369826 559286 369900 559314
rect 369826 559028 369854 559286
rect 379532 559042 379560 700538
rect 381188 700398 381216 703520
rect 390560 700528 390612 700534
rect 390560 700470 390612 700476
rect 381176 700392 381228 700398
rect 381176 700334 381228 700340
rect 390572 559042 390600 700470
rect 397472 700330 397500 703520
rect 413664 701010 413692 703520
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 429856 700942 429884 703520
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 446140 700874 446168 703520
rect 446128 700868 446180 700874
rect 446128 700810 446180 700816
rect 462332 700806 462360 703520
rect 462320 700800 462372 700806
rect 462320 700742 462372 700748
rect 478524 700738 478552 703520
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 511000 700602 511028 703520
rect 510988 700596 511040 700602
rect 510988 700538 511040 700544
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 401600 700460 401652 700466
rect 401600 700402 401652 700408
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 401612 559042 401640 700402
rect 559668 700398 559696 703520
rect 412640 700392 412692 700398
rect 412640 700334 412692 700340
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 412652 559042 412680 700334
rect 575860 700330 575888 703520
rect 423680 700324 423732 700330
rect 423680 700266 423732 700272
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 423692 559042 423720 700266
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 428464 683188 428516 683194
rect 428464 683130 428516 683136
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 379532 559014 380860 559042
rect 390572 559014 391860 559042
rect 401612 559014 402860 559042
rect 412652 559014 413840 559042
rect 423692 559014 424220 559042
rect 37832 545080 37884 545086
rect 37832 545022 37884 545028
rect 37844 544649 37872 545022
rect 37830 544640 37886 544649
rect 37830 544575 37886 544584
rect 37924 541680 37976 541686
rect 37924 541622 37976 541628
rect 37556 536784 37608 536790
rect 37556 536726 37608 536732
rect 37568 536217 37596 536726
rect 37554 536208 37610 536217
rect 37554 536143 37610 536152
rect 37832 527128 37884 527134
rect 37832 527070 37884 527076
rect 37844 526697 37872 527070
rect 37830 526688 37886 526697
rect 37830 526623 37886 526632
rect 37556 507816 37608 507822
rect 37556 507758 37608 507764
rect 37568 507521 37596 507758
rect 37554 507512 37610 507521
rect 37554 507447 37610 507456
rect 37936 498137 37964 541622
rect 428476 535401 428504 683130
rect 579618 630864 579674 630873
rect 579618 630799 579674 630808
rect 579632 630698 579660 630799
rect 428556 630692 428608 630698
rect 428556 630634 428608 630640
rect 579620 630692 579672 630698
rect 579620 630634 579672 630640
rect 428462 535392 428518 535401
rect 428462 535327 428518 535336
rect 428464 524476 428516 524482
rect 428464 524418 428516 524424
rect 38016 517472 38068 517478
rect 38016 517414 38068 517420
rect 38028 517177 38056 517414
rect 38014 517168 38070 517177
rect 38014 517103 38070 517112
rect 37922 498128 37978 498137
rect 37922 498063 37978 498072
rect 37832 488504 37884 488510
rect 37830 488472 37832 488481
rect 37884 488472 37886 488481
rect 37830 488407 37886 488416
rect 36542 478408 36598 478417
rect 36542 478343 36598 478352
rect 31024 474768 31076 474774
rect 31024 474710 31076 474716
rect 28264 422272 28316 422278
rect 28264 422214 28316 422220
rect 31036 383654 31064 474710
rect 37924 469192 37976 469198
rect 37924 469134 37976 469140
rect 37936 468897 37964 469134
rect 37922 468888 37978 468897
rect 37922 468823 37978 468832
rect 37464 459536 37516 459542
rect 37464 459478 37516 459484
rect 37476 459377 37504 459478
rect 37462 459368 37518 459377
rect 37462 459303 37518 459312
rect 37924 449880 37976 449886
rect 37922 449848 37924 449857
rect 37976 449848 37978 449857
rect 37922 449783 37978 449792
rect 37832 441584 37884 441590
rect 37832 441526 37884 441532
rect 37844 440881 37872 441526
rect 37830 440872 37886 440881
rect 37830 440807 37886 440816
rect 37832 431928 37884 431934
rect 37832 431870 37884 431876
rect 37844 431361 37872 431870
rect 37830 431352 37886 431361
rect 37830 431287 37886 431296
rect 37924 422272 37976 422278
rect 37924 422214 37976 422220
rect 37936 421841 37964 422214
rect 37922 421832 37978 421841
rect 37922 421767 37978 421776
rect 428476 419529 428504 524418
rect 428568 496777 428596 630634
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 428648 576904 428700 576910
rect 428648 576846 428700 576852
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 428554 496768 428610 496777
rect 428554 496703 428610 496712
rect 428556 487144 428608 487150
rect 428554 487112 428556 487121
rect 428608 487112 428610 487121
rect 428554 487047 428610 487056
rect 428556 477488 428608 477494
rect 428554 477456 428556 477465
rect 428608 477456 428610 477465
rect 428554 477391 428610 477400
rect 428556 470620 428608 470626
rect 428556 470562 428608 470568
rect 428462 419520 428518 419529
rect 428462 419455 428518 419464
rect 37648 412616 37700 412622
rect 37648 412558 37700 412564
rect 37660 412321 37688 412558
rect 37646 412312 37702 412321
rect 37646 412247 37702 412256
rect 37556 402960 37608 402966
rect 37556 402902 37608 402908
rect 37568 402529 37596 402902
rect 37554 402520 37610 402529
rect 37554 402455 37610 402464
rect 428464 400172 428516 400178
rect 428464 400114 428516 400120
rect 428476 399945 428504 400114
rect 428462 399936 428518 399945
rect 428462 399871 428518 399880
rect 37740 393304 37792 393310
rect 37740 393246 37792 393252
rect 37752 393145 37780 393246
rect 37738 393136 37794 393145
rect 37738 393071 37794 393080
rect 428464 390516 428516 390522
rect 428464 390458 428516 390464
rect 428476 390153 428504 390458
rect 428462 390144 428518 390153
rect 428462 390079 428518 390088
rect 31024 383648 31076 383654
rect 37464 383648 37516 383654
rect 31024 383590 31076 383596
rect 37462 383616 37464 383625
rect 37516 383616 37518 383625
rect 37462 383551 37518 383560
rect 428568 380633 428596 470562
rect 428660 458153 428688 576846
rect 580170 551168 580226 551177
rect 580170 551103 580226 551112
rect 580184 550662 580212 551103
rect 490564 550656 490616 550662
rect 490564 550598 490616 550604
rect 580172 550656 580224 550662
rect 580172 550598 580224 550604
rect 428740 545080 428792 545086
rect 428740 545022 428792 545028
rect 428752 544921 428780 545022
rect 428738 544912 428794 544921
rect 428738 544847 428794 544856
rect 428740 525768 428792 525774
rect 428738 525736 428740 525745
rect 428792 525736 428794 525745
rect 428738 525671 428794 525680
rect 428740 516112 428792 516118
rect 428738 516080 428740 516089
rect 428792 516080 428794 516089
rect 428738 516015 428794 516024
rect 428740 506456 428792 506462
rect 428738 506424 428740 506433
rect 428792 506424 428794 506433
rect 428738 506359 428794 506368
rect 428740 467832 428792 467838
rect 428738 467800 428740 467809
rect 428792 467800 428794 467809
rect 428738 467735 428794 467744
rect 428646 458144 428702 458153
rect 428646 458079 428702 458088
rect 429108 448520 429160 448526
rect 429108 448462 429160 448468
rect 429120 448225 429148 448462
rect 429106 448216 429162 448225
rect 429106 448151 429162 448160
rect 490576 438870 490604 550598
rect 580276 545086 580304 697167
rect 580354 670712 580410 670721
rect 580354 670647 580410 670656
rect 580264 545080 580316 545086
rect 580264 545022 580316 545028
rect 580262 537840 580318 537849
rect 580262 537775 580318 537784
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 428648 438864 428700 438870
rect 428648 438806 428700 438812
rect 490564 438864 490616 438870
rect 490564 438806 490616 438812
rect 428660 438705 428688 438806
rect 428646 438696 428702 438705
rect 428646 438631 428702 438640
rect 580078 431624 580134 431633
rect 580078 431559 580134 431568
rect 580092 430642 580120 431559
rect 428740 430636 428792 430642
rect 428740 430578 428792 430584
rect 580080 430636 580132 430642
rect 580080 430578 580132 430584
rect 428648 429140 428700 429146
rect 428648 429082 428700 429088
rect 428660 429049 428688 429082
rect 428646 429040 428702 429049
rect 428646 428975 428702 428984
rect 428752 422294 428780 430578
rect 580276 429146 580304 537775
rect 580368 525774 580396 670647
rect 580446 657384 580502 657393
rect 580446 657319 580502 657328
rect 580356 525768 580408 525774
rect 580356 525710 580408 525716
rect 580460 516118 580488 657319
rect 580538 644056 580594 644065
rect 580538 643991 580594 644000
rect 580448 516112 580500 516118
rect 580448 516054 580500 516060
rect 580354 511320 580410 511329
rect 580354 511255 580410 511264
rect 580264 429140 580316 429146
rect 580264 429082 580316 429088
rect 428660 422266 428780 422294
rect 428554 380624 428610 380633
rect 428554 380559 428610 380568
rect 37924 373992 37976 373998
rect 37922 373960 37924 373969
rect 37976 373960 37978 373969
rect 37922 373895 37978 373904
rect 428464 364404 428516 364410
rect 428464 364346 428516 364352
rect 37464 364336 37516 364342
rect 37464 364278 37516 364284
rect 37476 364177 37504 364278
rect 37462 364168 37518 364177
rect 37462 364103 37518 364112
rect 37556 354680 37608 354686
rect 37556 354622 37608 354628
rect 37568 354521 37596 354622
rect 37554 354512 37610 354521
rect 37554 354447 37610 354456
rect 26884 345024 26936 345030
rect 37648 345024 37700 345030
rect 26884 344966 26936 344972
rect 37646 344992 37648 345001
rect 37700 344992 37702 345001
rect 37646 344927 37702 344936
rect 37832 336728 37884 336734
rect 37832 336670 37884 336676
rect 37844 336025 37872 336670
rect 37830 336016 37886 336025
rect 37830 335951 37886 335960
rect 37556 327072 37608 327078
rect 37556 327014 37608 327020
rect 37568 326505 37596 327014
rect 37554 326496 37610 326505
rect 37554 326431 37610 326440
rect 24124 317416 24176 317422
rect 24124 317358 24176 317364
rect 37924 317416 37976 317422
rect 37924 317358 37976 317364
rect 37936 316985 37964 317358
rect 37922 316976 37978 316985
rect 37922 316911 37978 316920
rect 6184 307760 6236 307766
rect 6184 307702 6236 307708
rect 37372 307760 37424 307766
rect 37372 307702 37424 307708
rect 37384 307329 37412 307702
rect 37370 307320 37426 307329
rect 37370 307255 37426 307264
rect 428476 302841 428504 364346
rect 428556 361548 428608 361554
rect 428556 361490 428608 361496
rect 428568 361185 428596 361490
rect 428554 361176 428610 361185
rect 428554 361111 428610 361120
rect 428660 351393 428688 422266
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 428740 418192 428792 418198
rect 428740 418134 428792 418140
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 428646 351384 428702 351393
rect 428646 351319 428702 351328
rect 428752 341737 428780 418134
rect 580368 409834 580396 511255
rect 580552 506462 580580 643991
rect 580630 617536 580686 617545
rect 580630 617471 580686 617480
rect 580540 506456 580592 506462
rect 580540 506398 580592 506404
rect 580446 497992 580502 498001
rect 580446 497927 580502 497936
rect 428832 409828 428884 409834
rect 428832 409770 428884 409776
rect 580356 409828 580408 409834
rect 580356 409770 580408 409776
rect 428844 409465 428872 409770
rect 428830 409456 428886 409465
rect 428830 409391 428886 409400
rect 580262 404968 580318 404977
rect 580262 404903 580318 404912
rect 428832 371204 428884 371210
rect 428832 371146 428884 371152
rect 428844 370705 428872 371146
rect 428830 370696 428886 370705
rect 428830 370631 428886 370640
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 428738 341728 428794 341737
rect 428738 341663 428794 341672
rect 580276 332586 580304 404903
rect 580460 400178 580488 497927
rect 580644 487150 580672 617471
rect 580722 604208 580778 604217
rect 580722 604143 580778 604152
rect 580632 487144 580684 487150
rect 580632 487086 580684 487092
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580448 400172 580500 400178
rect 580448 400114 580500 400120
rect 580354 391776 580410 391785
rect 580354 391711 580410 391720
rect 428556 332580 428608 332586
rect 428556 332522 428608 332528
rect 580264 332580 580316 332586
rect 580264 332522 580316 332528
rect 428568 332081 428596 332522
rect 428554 332072 428610 332081
rect 428554 332007 428610 332016
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 324358 579660 325207
rect 428556 324352 428608 324358
rect 428556 324294 428608 324300
rect 579620 324352 579672 324358
rect 579620 324294 579672 324300
rect 428462 302832 428518 302841
rect 428462 302767 428518 302776
rect 37556 298104 37608 298110
rect 37556 298046 37608 298052
rect 37568 297673 37596 298046
rect 37554 297664 37610 297673
rect 37554 297599 37610 297608
rect 428464 292528 428516 292534
rect 428462 292496 428464 292505
rect 428516 292496 428518 292505
rect 428462 292431 428518 292440
rect 37740 288380 37792 288386
rect 37740 288322 37792 288328
rect 37752 288289 37780 288322
rect 37738 288280 37794 288289
rect 37738 288215 37794 288224
rect 4804 278724 4856 278730
rect 4804 278666 4856 278672
rect 37740 278724 37792 278730
rect 37740 278666 37792 278672
rect 37752 278497 37780 278666
rect 37738 278488 37794 278497
rect 37738 278423 37794 278432
rect 428568 273193 428596 324294
rect 580368 322930 580396 391711
rect 580552 390522 580580 484599
rect 580736 477494 580764 604143
rect 580814 591016 580870 591025
rect 580814 590951 580870 590960
rect 580724 477488 580776 477494
rect 580724 477430 580776 477436
rect 580828 470594 580856 590951
rect 580906 564360 580962 564369
rect 580906 564295 580962 564304
rect 580736 470566 580856 470594
rect 580736 467838 580764 470566
rect 580724 467832 580776 467838
rect 580724 467774 580776 467780
rect 580630 458144 580686 458153
rect 580630 458079 580686 458088
rect 580540 390516 580592 390522
rect 580540 390458 580592 390464
rect 580446 378448 580502 378457
rect 580446 378383 580502 378392
rect 428832 322924 428884 322930
rect 428832 322866 428884 322872
rect 580356 322924 580408 322930
rect 580356 322866 580408 322872
rect 428844 322289 428872 322866
rect 428830 322280 428886 322289
rect 428830 322215 428886 322224
rect 580460 313274 580488 378383
rect 580644 371210 580672 458079
rect 580920 448526 580948 564295
rect 580908 448520 580960 448526
rect 580908 448462 580960 448468
rect 580722 444816 580778 444825
rect 580722 444751 580778 444760
rect 580632 371204 580684 371210
rect 580632 371146 580684 371152
rect 580736 361554 580764 444751
rect 580724 361548 580776 361554
rect 580724 361490 580776 361496
rect 580538 351928 580594 351937
rect 580538 351863 580594 351872
rect 428740 313268 428792 313274
rect 428740 313210 428792 313216
rect 580448 313268 580500 313274
rect 580448 313210 580500 313216
rect 428752 312633 428780 313210
rect 428738 312624 428794 312633
rect 428738 312559 428794 312568
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 428648 311908 428700 311914
rect 428648 311850 428700 311856
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 428554 273184 428610 273193
rect 428554 273119 428610 273128
rect 428464 271924 428516 271930
rect 428464 271866 428516 271872
rect 37924 269068 37976 269074
rect 37924 269010 37976 269016
rect 37936 268977 37964 269010
rect 37922 268968 37978 268977
rect 37922 268903 37978 268912
rect 37372 259412 37424 259418
rect 37372 259354 37424 259360
rect 37384 258097 37412 259354
rect 37370 258088 37426 258097
rect 37370 258023 37426 258032
rect 37924 249756 37976 249762
rect 37924 249698 37976 249704
rect 37936 249665 37964 249698
rect 37922 249656 37978 249665
rect 37922 249591 37978 249600
rect 37370 240136 37426 240145
rect 3700 240100 3752 240106
rect 37370 240071 37372 240080
rect 3700 240042 3752 240048
rect 37424 240071 37426 240080
rect 37372 240042 37424 240048
rect 428476 234569 428504 271866
rect 428660 263537 428688 311850
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 429016 282872 429068 282878
rect 429014 282840 429016 282849
rect 429068 282840 429070 282849
rect 429014 282775 429070 282784
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579632 271930 579660 272167
rect 579620 271924 579672 271930
rect 579620 271866 579672 271872
rect 428646 263528 428702 263537
rect 428646 263463 428702 263472
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579632 258126 579660 258839
rect 428556 258120 428608 258126
rect 428556 258062 428608 258068
rect 579620 258120 579672 258126
rect 579620 258062 579672 258068
rect 428462 234560 428518 234569
rect 428462 234495 428518 234504
rect 428464 231872 428516 231878
rect 428464 231814 428516 231820
rect 37648 231804 37700 231810
rect 37648 231746 37700 231752
rect 37660 230625 37688 231746
rect 37646 230616 37702 230625
rect 37646 230551 37702 230560
rect 3608 222148 3660 222154
rect 3608 222090 3660 222096
rect 37740 222148 37792 222154
rect 37740 222090 37792 222096
rect 37752 221649 37780 222090
rect 37738 221640 37794 221649
rect 37738 221575 37794 221584
rect 3606 214976 3662 214985
rect 3606 214911 3662 214920
rect 3516 212492 3568 212498
rect 3516 212434 3568 212440
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3436 173874 3464 188799
rect 3528 183530 3556 201855
rect 3620 193186 3648 214911
rect 37832 212492 37884 212498
rect 37832 212434 37884 212440
rect 37844 212129 37872 212434
rect 37830 212120 37886 212129
rect 37830 212055 37886 212064
rect 428476 205601 428504 231814
rect 428568 224913 428596 258062
rect 580276 253910 580304 298687
rect 580552 292534 580580 351863
rect 580630 338600 580686 338609
rect 580630 338535 580686 338544
rect 580540 292528 580592 292534
rect 580540 292470 580592 292476
rect 580354 285424 580410 285433
rect 580354 285359 580410 285368
rect 428924 253904 428976 253910
rect 428922 253872 428924 253881
rect 580264 253904 580316 253910
rect 428976 253872 428978 253881
rect 580264 253846 580316 253852
rect 428922 253807 428978 253816
rect 579802 245576 579858 245585
rect 579802 245511 579858 245520
rect 579816 244322 579844 245511
rect 428740 244316 428792 244322
rect 428740 244258 428792 244264
rect 579804 244316 579856 244322
rect 579804 244258 579856 244264
rect 428648 244248 428700 244254
rect 428646 244216 428648 244225
rect 428700 244216 428702 244225
rect 428646 244151 428702 244160
rect 428752 238754 428780 244258
rect 580368 244254 580396 285359
rect 580644 282878 580672 338535
rect 580632 282872 580684 282878
rect 580632 282814 580684 282820
rect 580356 244248 580408 244254
rect 580356 244190 580408 244196
rect 428660 238726 428780 238754
rect 428554 224904 428610 224913
rect 428554 224839 428610 224848
rect 428556 218068 428608 218074
rect 428556 218010 428608 218016
rect 428462 205592 428518 205601
rect 428462 205527 428518 205536
rect 37740 202836 37792 202842
rect 37740 202778 37792 202784
rect 37752 202609 37780 202778
rect 37738 202600 37794 202609
rect 37738 202535 37794 202544
rect 428568 195945 428596 218010
rect 428660 215257 428688 238726
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 428646 215248 428702 215257
rect 428646 215183 428702 215192
rect 580170 205728 580226 205737
rect 428648 205692 428700 205698
rect 580170 205663 580172 205672
rect 428648 205634 428700 205640
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 428554 195936 428610 195945
rect 428554 195871 428610 195880
rect 3608 193180 3660 193186
rect 3608 193122 3660 193128
rect 37740 193180 37792 193186
rect 37740 193122 37792 193128
rect 37752 192953 37780 193122
rect 37738 192944 37794 192953
rect 37738 192879 37794 192888
rect 428464 191888 428516 191894
rect 428464 191830 428516 191836
rect 3516 183524 3568 183530
rect 3516 183466 3568 183472
rect 37924 183524 37976 183530
rect 37924 183466 37976 183472
rect 37936 183433 37964 183466
rect 37922 183424 37978 183433
rect 37922 183359 37978 183368
rect 428476 176633 428504 191830
rect 428660 186289 428688 205634
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 428646 186280 428702 186289
rect 428646 186215 428702 186224
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 428556 178084 428608 178090
rect 428556 178026 428608 178032
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 428462 176624 428518 176633
rect 428462 176559 428518 176568
rect 3514 175944 3570 175953
rect 3514 175879 3570 175888
rect 3424 173868 3476 173874
rect 3424 173810 3476 173816
rect 3528 164218 3556 175879
rect 37740 173868 37792 173874
rect 37740 173810 37792 173816
rect 37752 173641 37780 173810
rect 37738 173632 37794 173641
rect 37738 173567 37794 173576
rect 428568 166841 428596 178026
rect 428554 166832 428610 166841
rect 428554 166767 428610 166776
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 428464 165640 428516 165646
rect 428464 165582 428516 165588
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 3516 164212 3568 164218
rect 3516 164154 3568 164160
rect 37924 164212 37976 164218
rect 37924 164154 37976 164160
rect 37936 164121 37964 164154
rect 37922 164112 37978 164121
rect 37922 164047 37978 164056
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3436 154562 3464 162823
rect 428476 157185 428504 165582
rect 428462 157176 428518 157185
rect 428462 157111 428518 157120
rect 3424 154556 3476 154562
rect 3424 154498 3476 154504
rect 37648 154556 37700 154562
rect 37648 154498 37700 154504
rect 37660 154329 37688 154498
rect 37646 154320 37702 154329
rect 37646 154255 37702 154264
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 429108 151836 429160 151842
rect 429108 151778 429160 151784
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 144906 3372 149767
rect 429120 147393 429148 151778
rect 429106 147384 429162 147393
rect 429106 147319 429162 147328
rect 3332 144900 3384 144906
rect 3332 144842 3384 144848
rect 37924 144900 37976 144906
rect 37924 144842 37976 144848
rect 37936 144809 37964 144842
rect 37922 144800 37978 144809
rect 37922 144735 37978 144744
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 428832 138032 428884 138038
rect 428832 137974 428884 137980
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 428844 137601 428872 137974
rect 428830 137592 428886 137601
rect 428830 137527 428886 137536
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3436 136610 3464 136711
rect 3424 136604 3476 136610
rect 3424 136546 3476 136552
rect 37556 136604 37608 136610
rect 37556 136546 37608 136552
rect 37568 135833 37596 136546
rect 37554 135824 37610 135833
rect 37554 135759 37610 135768
rect 428922 127120 428978 127129
rect 428922 127055 428978 127064
rect 428936 126954 428964 127055
rect 428924 126948 428976 126954
rect 428924 126890 428976 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 37738 125760 37794 125769
rect 37738 125695 37794 125704
rect 37752 124166 37780 125695
rect 3424 124160 3476 124166
rect 3424 124102 3476 124108
rect 37740 124160 37792 124166
rect 37740 124102 37792 124108
rect 3436 123729 3464 124102
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 428462 117328 428518 117337
rect 428462 117263 428518 117272
rect 37922 115968 37978 115977
rect 37922 115903 37978 115912
rect 37936 111790 37964 115903
rect 428476 113150 428504 117263
rect 428464 113144 428516 113150
rect 428464 113086 428516 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 37924 111784 37976 111790
rect 37924 111726 37976 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 428462 107672 428518 107681
rect 428462 107607 428518 107616
rect 37922 106312 37978 106321
rect 37922 106247 37978 106256
rect 37936 97986 37964 106247
rect 428476 100706 428504 107607
rect 428464 100700 428516 100706
rect 428464 100642 428516 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 428554 98016 428610 98025
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 37924 97980 37976 97986
rect 428554 97951 428610 97960
rect 37924 97922 37976 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 38014 96656 38070 96665
rect 38014 96591 38070 96600
rect 37922 87000 37978 87009
rect 37922 86935 37978 86944
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 37936 71738 37964 86935
rect 38028 85542 38056 96591
rect 428462 88360 428518 88369
rect 428462 88295 428518 88304
rect 38016 85536 38068 85542
rect 38016 85478 38068 85484
rect 38014 77480 38070 77489
rect 38014 77415 38070 77424
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 37924 71732 37976 71738
rect 37924 71674 37976 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 37922 67960 37978 67969
rect 37922 67895 37978 67904
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 37936 45558 37964 67895
rect 38028 59362 38056 77415
rect 428476 73166 428504 88295
rect 428568 86970 428596 97951
rect 428556 86964 428608 86970
rect 428556 86906 428608 86912
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 428554 78704 428610 78713
rect 428554 78639 428610 78648
rect 428464 73160 428516 73166
rect 428464 73102 428516 73108
rect 428462 69184 428518 69193
rect 428462 69119 428518 69128
rect 38016 59356 38068 59362
rect 38016 59298 38068 59304
rect 38106 58440 38162 58449
rect 38106 58375 38162 58384
rect 38014 49328 38070 49337
rect 38014 49263 38070 49272
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 37924 45552 37976 45558
rect 3476 45520 3478 45529
rect 37924 45494 37976 45500
rect 3422 45455 3478 45464
rect 37922 40216 37978 40225
rect 37922 40151 37978 40160
rect 10324 37936 10376 37942
rect 10324 37878 10376 37884
rect 4804 36644 4856 36650
rect 4804 36586 4856 36592
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 2780 28280 2832 28286
rect 2780 28222 2832 28228
rect 2792 16574 2820 28222
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2792 16546 3648 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 480 1716 2994
rect 2884 480 2912 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 3058 4016 8910
rect 4816 3534 4844 36586
rect 6920 35216 6972 35222
rect 6920 35158 6972 35164
rect 6932 16574 6960 35158
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8312 16574 8340 17206
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 5276 480 5304 3295
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9968 480 9996 3538
rect 10336 3466 10364 37878
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 11060 33788 11112 33794
rect 11060 33730 11112 33736
rect 11072 16574 11100 33730
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 11072 16546 11928 16574
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 14476 3534 14504 26862
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13556 480 13584 3470
rect 14752 480 14780 4082
rect 15856 3602 15884 29582
rect 17040 10328 17092 10334
rect 17040 10270 17092 10276
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15948 480 15976 3470
rect 17052 480 17080 10270
rect 17236 4146 17264 36518
rect 35900 32428 35952 32434
rect 35900 32370 35952 32376
rect 20720 31204 20772 31210
rect 20720 31146 20772 31152
rect 17960 25560 18012 25566
rect 17960 25502 18012 25508
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 25502
rect 20732 16574 20760 31146
rect 33140 29708 33192 29714
rect 33140 29650 33192 29656
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22112 16574 22140 24074
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27632 16574 27660 21422
rect 33152 16574 33180 29650
rect 34520 22840 34572 22846
rect 34520 22782 34572 22788
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 27632 16546 27752 16574
rect 33152 16546 33640 16574
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19444 480 19472 3674
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20640 480 20668 3538
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 26516 7608 26568 7614
rect 26516 7550 26568 7556
rect 24216 3800 24268 3806
rect 24216 3742 24268 3748
rect 24228 480 24256 3742
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25332 480 25360 3606
rect 26528 480 26556 7550
rect 27724 480 27752 16546
rect 30840 14544 30892 14550
rect 30840 14486 30892 14492
rect 30104 13116 30156 13122
rect 30104 13058 30156 13064
rect 28908 3868 28960 3874
rect 28908 3810 28960 3816
rect 28920 480 28948 3810
rect 30116 480 30144 13058
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 14486
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32416 480 32444 3878
rect 33612 480 33640 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 22782
rect 35912 16574 35940 32370
rect 35912 16546 36768 16574
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 36004 480 36032 3946
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 37832 11824 37884 11830
rect 37832 11766 37884 11772
rect 37844 3482 37872 11766
rect 37936 6866 37964 40151
rect 38028 20670 38056 49263
rect 38120 33114 38148 58375
rect 428476 46918 428504 69119
rect 428568 60722 428596 78639
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 428556 60716 428608 60722
rect 428556 60658 428608 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 428646 59392 428702 59401
rect 428646 59327 428702 59336
rect 428554 49056 428610 49065
rect 428554 48991 428610 49000
rect 428464 46912 428516 46918
rect 428464 46854 428516 46860
rect 67652 40174 68416 40202
rect 42812 40140 43484 40168
rect 40144 40034 40400 40062
rect 40512 40035 40760 40063
rect 41432 40035 41520 40063
rect 41984 40035 42300 40063
rect 39304 38004 39356 38010
rect 39304 37946 39356 37952
rect 38108 33108 38160 33114
rect 38108 33050 38160 33056
rect 38016 20664 38068 20670
rect 38016 20606 38068 20612
rect 37924 6860 37976 6866
rect 37924 6802 37976 6808
rect 39316 4826 39344 37946
rect 40144 8974 40172 40034
rect 40512 38010 40540 40035
rect 40500 38004 40552 38010
rect 40500 37946 40552 37952
rect 41328 38004 41380 38010
rect 41328 37946 41380 37952
rect 41340 35222 41368 37946
rect 41432 36650 41460 40035
rect 41984 38010 42012 40035
rect 41972 38004 42024 38010
rect 41972 37946 42024 37952
rect 41420 36644 41472 36650
rect 41420 36586 41472 36592
rect 41328 35216 41380 35222
rect 41328 35158 41380 35164
rect 41880 10396 41932 10402
rect 41880 10338 41932 10344
rect 40132 8968 40184 8974
rect 40132 8910 40184 8916
rect 39304 4820 39356 4826
rect 39304 4762 39356 4768
rect 40684 4616 40736 4622
rect 40684 4558 40736 4564
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 37844 3454 38424 3482
rect 38396 480 38424 3454
rect 39592 480 39620 4014
rect 40696 480 40724 4558
rect 41892 480 41920 10338
rect 42812 10334 42840 40140
rect 43456 40066 43484 40140
rect 42904 40035 43080 40063
rect 43456 40038 43860 40066
rect 44284 40035 44640 40063
rect 45112 40035 45440 40063
rect 45756 40035 46220 40063
rect 42904 33794 42932 40035
rect 44180 38004 44232 38010
rect 44180 37946 44232 37952
rect 42892 33788 42944 33794
rect 42892 33730 42944 33736
rect 42800 10328 42852 10334
rect 42800 10270 42852 10276
rect 44192 7614 44220 37946
rect 44284 31210 44312 40035
rect 45112 38010 45140 40035
rect 45100 38004 45152 38010
rect 45100 37946 45152 37952
rect 44272 31204 44324 31210
rect 44272 31146 44324 31152
rect 44272 31068 44324 31074
rect 44272 31010 44324 31016
rect 44284 16574 44312 31010
rect 45756 26234 45784 40035
rect 46986 39794 47014 40049
rect 46952 39766 47014 39794
rect 47412 40035 47780 40063
rect 48332 40035 48560 40063
rect 48976 40035 49340 40063
rect 49804 40035 50120 40063
rect 50632 40035 50920 40063
rect 51276 40035 51700 40063
rect 52480 40035 52592 40063
rect 46204 38276 46256 38282
rect 46204 38218 46256 38224
rect 45572 26206 45784 26234
rect 44284 16546 45048 16574
rect 44180 7608 44232 7614
rect 44180 7550 44232 7556
rect 44272 5568 44324 5574
rect 44272 5510 44324 5516
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 43088 480 43116 4082
rect 44284 480 44312 5510
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 45572 13122 45600 26206
rect 45560 13116 45612 13122
rect 45560 13058 45612 13064
rect 46216 5574 46244 38218
rect 46952 29714 46980 39766
rect 47412 32434 47440 40035
rect 48332 38350 48360 40035
rect 47584 38344 47636 38350
rect 47584 38286 47636 38292
rect 48320 38344 48372 38350
rect 48320 38286 48372 38292
rect 47400 32428 47452 32434
rect 47400 32370 47452 32376
rect 46940 29708 46992 29714
rect 46940 29650 46992 29656
rect 46204 5568 46256 5574
rect 46204 5510 46256 5516
rect 47596 4622 47624 38286
rect 48976 38282 49004 40035
rect 48964 38276 49016 38282
rect 48964 38218 49016 38224
rect 49700 38004 49752 38010
rect 49700 37946 49752 37952
rect 48320 18692 48372 18698
rect 48320 18634 48372 18640
rect 48332 16574 48360 18634
rect 48332 16546 48544 16574
rect 47584 4616 47636 4622
rect 47584 4558 47636 4564
rect 47860 4208 47912 4214
rect 47860 4150 47912 4156
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 46676 480 46704 3334
rect 47872 480 47900 4150
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 49712 4282 49740 37946
rect 49700 4276 49752 4282
rect 49700 4218 49752 4224
rect 49804 4214 49832 40035
rect 50632 38010 50660 40035
rect 50620 38004 50672 38010
rect 50620 37946 50672 37952
rect 49884 32428 49936 32434
rect 49884 32370 49936 32376
rect 49896 16574 49924 32370
rect 51276 26234 51304 40035
rect 52460 38004 52512 38010
rect 52460 37946 52512 37952
rect 51092 26206 51304 26234
rect 49896 16546 50200 16574
rect 49792 4208 49844 4214
rect 49792 4150 49844 4156
rect 50172 480 50200 16546
rect 51092 4214 51120 26206
rect 52472 4826 52500 37946
rect 52564 6186 52592 40035
rect 52932 40035 53240 40063
rect 53852 40035 54020 40063
rect 54404 40035 54800 40063
rect 55580 40035 55904 40063
rect 56360 40035 56548 40063
rect 52932 38010 52960 40035
rect 52920 38004 52972 38010
rect 52920 37946 52972 37952
rect 52644 20052 52696 20058
rect 52644 19994 52696 20000
rect 52552 6180 52604 6186
rect 52552 6122 52604 6128
rect 52460 4820 52512 4826
rect 52460 4762 52512 4768
rect 51356 4276 51408 4282
rect 51356 4218 51408 4224
rect 51080 4208 51132 4214
rect 51080 4150 51132 4156
rect 51368 480 51396 4218
rect 52656 1306 52684 19994
rect 53288 13116 53340 13122
rect 53288 13058 53340 13064
rect 52564 1278 52684 1306
rect 52564 480 52592 1278
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 13058
rect 53852 7682 53880 40035
rect 54404 26234 54432 40035
rect 55876 38418 55904 40035
rect 55864 38412 55916 38418
rect 55864 38354 55916 38360
rect 56520 36650 56548 40035
rect 56796 40035 57140 40063
rect 57624 40035 57920 40063
rect 58268 40035 58700 40063
rect 59480 40035 59768 40063
rect 56600 38004 56652 38010
rect 56600 37946 56652 37952
rect 56508 36644 56560 36650
rect 56508 36586 56560 36592
rect 55220 33788 55272 33794
rect 55220 33730 55272 33736
rect 53944 26206 54432 26234
rect 53944 9042 53972 26206
rect 55232 16574 55260 33730
rect 55232 16546 56088 16574
rect 53932 9036 53984 9042
rect 53932 8978 53984 8984
rect 53840 7676 53892 7682
rect 53840 7618 53892 7624
rect 54944 4208 54996 4214
rect 54944 4150 54996 4156
rect 54956 480 54984 4150
rect 56060 480 56088 16546
rect 56612 5030 56640 37946
rect 56796 26234 56824 40035
rect 57624 38010 57652 40035
rect 57612 38004 57664 38010
rect 57612 37946 57664 37952
rect 58268 26234 58296 40035
rect 58624 38412 58676 38418
rect 58624 38354 58676 38360
rect 56704 26206 56824 26234
rect 57992 26206 58296 26234
rect 56704 5098 56732 26206
rect 56784 21412 56836 21418
rect 56784 21354 56836 21360
rect 56692 5092 56744 5098
rect 56692 5034 56744 5040
rect 56600 5024 56652 5030
rect 56600 4966 56652 4972
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 21354
rect 57992 4962 58020 26206
rect 58636 6254 58664 38354
rect 59740 38078 59768 40035
rect 59832 40035 60260 40063
rect 60752 40035 61060 40063
rect 61396 40035 61840 40063
rect 62224 40035 62620 40063
rect 63144 40035 63400 40063
rect 63788 40035 64180 40063
rect 59728 38072 59780 38078
rect 59728 38014 59780 38020
rect 59832 26234 59860 40035
rect 59372 26206 59860 26234
rect 59372 15910 59400 26206
rect 59360 15904 59412 15910
rect 59360 15846 59412 15852
rect 60752 10334 60780 40035
rect 61396 26234 61424 40035
rect 62120 38004 62172 38010
rect 62120 37946 62172 37952
rect 60844 26206 61424 26234
rect 60844 11762 60872 26206
rect 60924 18624 60976 18630
rect 60924 18566 60976 18572
rect 60832 11756 60884 11762
rect 60832 11698 60884 11704
rect 60740 10328 60792 10334
rect 60740 10270 60792 10276
rect 59636 7608 59688 7614
rect 59636 7550 59688 7556
rect 58624 6248 58676 6254
rect 58624 6190 58676 6196
rect 58440 6180 58492 6186
rect 58440 6122 58492 6128
rect 57980 4956 58032 4962
rect 57980 4898 58032 4904
rect 58452 480 58480 6122
rect 59648 480 59676 7550
rect 60936 6914 60964 18566
rect 60844 6886 60964 6914
rect 60844 480 60872 6886
rect 62132 4826 62160 37946
rect 62224 4894 62252 40035
rect 63144 38010 63172 40035
rect 63132 38004 63184 38010
rect 63132 37946 63184 37952
rect 63788 26234 63816 40035
rect 64946 39794 64974 40049
rect 65444 40035 65740 40063
rect 66520 40035 66852 40063
rect 64946 39766 65012 39794
rect 64880 38004 64932 38010
rect 64880 37946 64932 37952
rect 63512 26206 63816 26234
rect 63512 13190 63540 26206
rect 63592 22772 63644 22778
rect 63592 22714 63644 22720
rect 63604 16574 63632 22714
rect 63604 16546 64368 16574
rect 63500 13184 63552 13190
rect 63500 13126 63552 13132
rect 63224 8968 63276 8974
rect 63224 8910 63276 8916
rect 62212 4888 62264 4894
rect 62212 4830 62264 4836
rect 62028 4820 62080 4826
rect 62028 4762 62080 4768
rect 62120 4820 62172 4826
rect 62120 4762 62172 4768
rect 62040 480 62068 4762
rect 63236 480 63264 8910
rect 64340 480 64368 16546
rect 64892 6186 64920 37946
rect 64984 14482 65012 39766
rect 65444 38010 65472 40035
rect 66824 38146 66852 40035
rect 66916 40035 67300 40063
rect 66812 38140 66864 38146
rect 66812 38082 66864 38088
rect 65432 38004 65484 38010
rect 65432 37946 65484 37952
rect 66916 28286 66944 40035
rect 66904 28280 66956 28286
rect 66904 28222 66956 28228
rect 67652 26926 67680 40174
rect 68388 40066 68416 40174
rect 82832 40174 83320 40202
rect 67744 40035 68080 40063
rect 68388 40038 68860 40066
rect 69216 40035 69640 40063
rect 70400 40035 70532 40063
rect 67640 26920 67692 26926
rect 67640 26862 67692 26868
rect 66260 17332 66312 17338
rect 66260 17274 66312 17280
rect 66272 16574 66300 17274
rect 67744 17270 67772 40035
rect 68928 38140 68980 38146
rect 68928 38082 68980 38088
rect 68940 35222 68968 38082
rect 68928 35216 68980 35222
rect 68928 35158 68980 35164
rect 67824 27056 67876 27062
rect 67824 26998 67876 27004
rect 67732 17264 67784 17270
rect 67732 17206 67784 17212
rect 67836 16574 67864 26998
rect 69216 26234 69244 40035
rect 69664 38072 69716 38078
rect 69664 38014 69716 38020
rect 69032 26206 69244 26234
rect 69032 25566 69060 26206
rect 69020 25560 69072 25566
rect 69020 25502 69072 25508
rect 66272 16546 66760 16574
rect 67836 16546 67956 16574
rect 64972 14476 65024 14482
rect 64972 14418 65024 14424
rect 65524 7676 65576 7682
rect 65524 7618 65576 7624
rect 64880 6180 64932 6186
rect 64880 6122 64932 6128
rect 65536 480 65564 7618
rect 66732 480 66760 16546
rect 67928 480 67956 16546
rect 69112 9036 69164 9042
rect 69112 8978 69164 8984
rect 69124 480 69152 8978
rect 69676 7682 69704 38014
rect 70400 38004 70452 38010
rect 70400 37946 70452 37952
rect 70412 21486 70440 37946
rect 70504 24138 70532 40035
rect 70872 40035 71200 40063
rect 71792 40035 71980 40063
rect 72344 40035 72760 40063
rect 73264 40035 73540 40063
rect 74000 40035 74320 40063
rect 74644 40035 75100 40063
rect 75564 40035 75880 40063
rect 76300 40035 76680 40063
rect 77312 40035 77440 40063
rect 77864 40035 78220 40063
rect 78692 40035 79000 40063
rect 79428 40035 79780 40063
rect 80164 40035 80560 40063
rect 80992 40035 81340 40063
rect 81728 40035 82140 40063
rect 70872 38010 70900 40035
rect 70860 38004 70912 38010
rect 70860 37946 70912 37952
rect 71044 38004 71096 38010
rect 71044 37946 71096 37952
rect 70584 24200 70636 24206
rect 70584 24142 70636 24148
rect 70492 24132 70544 24138
rect 70492 24074 70544 24080
rect 70400 21480 70452 21486
rect 70400 21422 70452 21428
rect 70308 9036 70360 9042
rect 70308 8978 70360 8984
rect 69664 7676 69716 7682
rect 69664 7618 69716 7624
rect 70320 480 70348 8978
rect 70596 6914 70624 24142
rect 71056 11830 71084 37946
rect 71792 14550 71820 40035
rect 72344 26234 72372 40035
rect 72424 38616 72476 38622
rect 72424 38558 72476 38564
rect 71884 26206 72372 26234
rect 71884 22846 71912 26206
rect 71872 22840 71924 22846
rect 71872 22782 71924 22788
rect 71780 14544 71832 14550
rect 71780 14486 71832 14492
rect 71044 11824 71096 11830
rect 71044 11766 71096 11772
rect 72436 10402 72464 38558
rect 73264 38010 73292 40035
rect 74000 38622 74028 40035
rect 73988 38616 74040 38622
rect 73988 38558 74040 38564
rect 73252 38004 73304 38010
rect 73252 37946 73304 37952
rect 74540 38004 74592 38010
rect 74540 37946 74592 37952
rect 74552 18698 74580 37946
rect 74644 31074 74672 40035
rect 75564 38010 75592 40035
rect 76300 39930 76328 40035
rect 76024 39902 76328 39930
rect 75920 38208 75972 38214
rect 75920 38150 75972 38156
rect 75552 38004 75604 38010
rect 75552 37946 75604 37952
rect 75184 37868 75236 37874
rect 75184 37810 75236 37816
rect 74632 31068 74684 31074
rect 74632 31010 74684 31016
rect 74632 19984 74684 19990
rect 74632 19926 74684 19932
rect 74540 18692 74592 18698
rect 74540 18634 74592 18640
rect 74644 16574 74672 19926
rect 74644 16546 75040 16574
rect 72424 10396 72476 10402
rect 72424 10338 72476 10344
rect 70596 6886 71544 6914
rect 71516 480 71544 6886
rect 72608 6248 72660 6254
rect 72608 6190 72660 6196
rect 73804 6248 73856 6254
rect 73804 6190 73856 6196
rect 72620 480 72648 6190
rect 73816 480 73844 6190
rect 75012 480 75040 16546
rect 75196 7614 75224 37810
rect 75932 33794 75960 38150
rect 75920 33788 75972 33794
rect 75920 33730 75972 33736
rect 76024 31210 76052 39902
rect 77312 38214 77340 40035
rect 77300 38208 77352 38214
rect 77300 38150 77352 38156
rect 77864 37874 77892 40035
rect 77852 37868 77904 37874
rect 77852 37810 77904 37816
rect 76104 36644 76156 36650
rect 76104 36586 76156 36592
rect 76012 31204 76064 31210
rect 76012 31146 76064 31152
rect 76116 31090 76144 36586
rect 75932 31062 76144 31090
rect 75184 7608 75236 7614
rect 75184 7550 75236 7556
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 31062
rect 76012 31000 76064 31006
rect 76012 30942 76064 30948
rect 76024 20058 76052 30942
rect 77300 25560 77352 25566
rect 77300 25502 77352 25508
rect 76012 20052 76064 20058
rect 76012 19994 76064 20000
rect 77312 16574 77340 25502
rect 77312 16546 78168 16574
rect 77392 7268 77444 7274
rect 77392 7210 77444 7216
rect 77404 480 77432 7210
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78692 8974 78720 40035
rect 79428 26234 79456 40035
rect 80060 38004 80112 38010
rect 80060 37946 80112 37952
rect 78784 26206 79456 26234
rect 78784 17338 78812 26206
rect 78772 17332 78824 17338
rect 78772 17274 78824 17280
rect 78680 8968 78732 8974
rect 78680 8910 78732 8916
rect 80072 6254 80100 37946
rect 80164 9042 80192 40035
rect 80992 38010 81020 40035
rect 80980 38004 81032 38010
rect 80980 37946 81032 37952
rect 81728 26234 81756 40035
rect 81452 26206 81756 26234
rect 80152 9036 80204 9042
rect 80152 8978 80204 8984
rect 80888 8764 80940 8770
rect 80888 8706 80940 8712
rect 80060 6248 80112 6254
rect 80060 6190 80112 6196
rect 79692 5092 79744 5098
rect 79692 5034 79744 5040
rect 79704 480 79732 5034
rect 80900 480 80928 8706
rect 81452 7274 81480 26206
rect 81624 15972 81676 15978
rect 81624 15914 81676 15920
rect 81440 7268 81492 7274
rect 81440 7210 81492 7216
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 15914
rect 82832 4350 82860 40174
rect 83292 40066 83320 40174
rect 100772 40174 101260 40202
rect 82920 40035 82952 40063
rect 83292 40038 83700 40066
rect 84460 40035 84792 40063
rect 82924 8770 82952 40035
rect 84764 38078 84792 40035
rect 84856 40035 85240 40063
rect 85684 40035 86020 40063
rect 86512 40035 86820 40063
rect 87156 40035 87600 40063
rect 88380 40035 88472 40063
rect 84752 38072 84804 38078
rect 84752 38014 84804 38020
rect 84856 26234 84884 40035
rect 85580 38004 85632 38010
rect 85580 37946 85632 37952
rect 84212 26206 84884 26234
rect 82912 8764 82964 8770
rect 82912 8706 82964 8712
rect 84212 5574 84240 26206
rect 85592 7750 85620 37946
rect 85684 16574 85712 40035
rect 86512 38010 86540 40035
rect 86960 38072 87012 38078
rect 86960 38014 87012 38020
rect 86500 38004 86552 38010
rect 86500 37946 86552 37952
rect 85684 16546 85804 16574
rect 85672 11824 85724 11830
rect 85672 11766 85724 11772
rect 85580 7744 85632 7750
rect 85580 7686 85632 7692
rect 84200 5568 84252 5574
rect 84200 5510 84252 5516
rect 83280 5024 83332 5030
rect 83280 4966 83332 4972
rect 82820 4344 82872 4350
rect 82820 4286 82872 4292
rect 83292 480 83320 4966
rect 84476 4344 84528 4350
rect 84476 4286 84528 4292
rect 84488 480 84516 4286
rect 85684 480 85712 11766
rect 85776 9110 85804 16546
rect 85764 9104 85816 9110
rect 85764 9046 85816 9052
rect 86972 6914 87000 38014
rect 87156 26234 87184 40035
rect 88340 38004 88392 38010
rect 88340 37946 88392 37952
rect 87064 26206 87184 26234
rect 87064 9042 87092 26206
rect 87052 9036 87104 9042
rect 87052 8978 87104 8984
rect 88352 7614 88380 37946
rect 88444 17270 88472 40035
rect 88904 40035 89160 40063
rect 89732 40035 89940 40063
rect 90700 40035 91048 40063
rect 91480 40035 91784 40063
rect 92280 40035 92428 40063
rect 88904 38010 88932 40035
rect 88892 38004 88944 38010
rect 88892 37946 88944 37952
rect 88432 17264 88484 17270
rect 88432 17206 88484 17212
rect 89732 10402 89760 40035
rect 91020 38078 91048 40035
rect 91008 38072 91060 38078
rect 91008 38014 91060 38020
rect 91756 38010 91784 40035
rect 91744 38004 91796 38010
rect 91744 37946 91796 37952
rect 92400 36650 92428 40035
rect 92676 40035 93060 40063
rect 93840 40038 93992 40066
rect 92388 36644 92440 36650
rect 92388 36586 92440 36592
rect 92676 29646 92704 40035
rect 93124 38072 93176 38078
rect 93124 38014 93176 38020
rect 92664 29640 92716 29646
rect 92664 29582 92716 29588
rect 89720 10396 89772 10402
rect 89720 10338 89772 10344
rect 93136 8974 93164 38014
rect 93964 36582 93992 40038
rect 94148 40035 94620 40063
rect 95252 40035 95400 40063
rect 95804 40035 96180 40063
rect 96632 40035 96960 40063
rect 97368 40035 97760 40063
rect 98104 40035 98520 40063
rect 99024 40035 99300 40063
rect 99668 40035 100080 40063
rect 93952 36576 94004 36582
rect 93952 36518 94004 36524
rect 94148 26234 94176 40035
rect 94056 26206 94176 26234
rect 93952 15904 94004 15910
rect 93952 15846 94004 15852
rect 93124 8968 93176 8974
rect 93124 8910 93176 8916
rect 90364 7676 90416 7682
rect 90364 7618 90416 7624
rect 88340 7608 88392 7614
rect 88340 7550 88392 7556
rect 86972 6886 87552 6914
rect 86868 4956 86920 4962
rect 86868 4898 86920 4904
rect 86880 480 86908 4898
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 6886
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 89180 480 89208 3266
rect 90376 480 90404 7618
rect 91560 5568 91612 5574
rect 91560 5510 91612 5516
rect 91572 480 91600 5510
rect 92756 3256 92808 3262
rect 92756 3198 92808 3204
rect 92768 480 92796 3198
rect 93964 480 93992 15846
rect 94056 3738 94084 26206
rect 95148 9104 95200 9110
rect 95148 9046 95200 9052
rect 94044 3732 94096 3738
rect 94044 3674 94096 3680
rect 95160 480 95188 9046
rect 95252 3806 95280 40035
rect 95804 26234 95832 40035
rect 95344 26206 95832 26234
rect 95344 3874 95372 26206
rect 96632 3942 96660 40035
rect 97368 26234 97396 40035
rect 98000 38072 98052 38078
rect 98000 38014 98052 38020
rect 96724 26206 97396 26234
rect 96724 4010 96752 26206
rect 97448 10328 97500 10334
rect 97448 10270 97500 10276
rect 96712 4004 96764 4010
rect 96712 3946 96764 3952
rect 96620 3936 96672 3942
rect 96620 3878 96672 3884
rect 95332 3868 95384 3874
rect 95332 3810 95384 3816
rect 95240 3800 95292 3806
rect 95240 3742 95292 3748
rect 96252 3732 96304 3738
rect 96252 3674 96304 3680
rect 96264 480 96292 3674
rect 97460 480 97488 10270
rect 98012 4146 98040 38014
rect 98000 4140 98052 4146
rect 98000 4082 98052 4088
rect 98104 4078 98132 40035
rect 99024 38078 99052 40035
rect 99012 38072 99064 38078
rect 99012 38014 99064 38020
rect 99668 26234 99696 40035
rect 99392 26206 99696 26234
rect 98644 7744 98696 7750
rect 98644 7686 98696 7692
rect 98092 4072 98144 4078
rect 98092 4014 98144 4020
rect 98656 480 98684 7686
rect 99392 3398 99420 26206
rect 100772 13122 100800 40174
rect 101232 40066 101260 40174
rect 107672 40174 108344 40202
rect 100860 40035 100892 40063
rect 101232 40038 101640 40066
rect 100864 32434 100892 40035
rect 102152 40035 102420 40063
rect 102796 40035 103200 40063
rect 103532 40035 103980 40063
rect 104360 40035 104760 40063
rect 105188 40035 105540 40063
rect 102152 38078 102180 40035
rect 101404 38072 101456 38078
rect 101404 38014 101456 38020
rect 102140 38072 102192 38078
rect 102140 38014 102192 38020
rect 100852 32428 100904 32434
rect 100852 32370 100904 32376
rect 101416 21418 101444 38014
rect 102796 26234 102824 40035
rect 102244 26206 102824 26234
rect 101404 21412 101456 21418
rect 101404 21354 101456 21360
rect 102244 18630 102272 26206
rect 103532 22778 103560 40035
rect 104360 38706 104388 40035
rect 104084 38678 104388 38706
rect 104084 27062 104112 38678
rect 104164 38004 104216 38010
rect 104164 37946 104216 37952
rect 104072 27056 104124 27062
rect 104072 26998 104124 27004
rect 103520 22772 103572 22778
rect 103520 22714 103572 22720
rect 104176 19990 104204 37946
rect 105188 26234 105216 40035
rect 105544 38072 105596 38078
rect 105544 38014 105596 38020
rect 104912 26206 105216 26234
rect 104912 24206 104940 26206
rect 104900 24200 104952 24206
rect 104900 24142 104952 24148
rect 104164 19984 104216 19990
rect 104164 19926 104216 19932
rect 102232 18624 102284 18630
rect 102232 18566 102284 18572
rect 104900 17264 104952 17270
rect 104900 17206 104952 17212
rect 100760 13116 100812 13122
rect 100760 13058 100812 13064
rect 100760 11756 100812 11762
rect 100760 11698 100812 11704
rect 99840 3800 99892 3806
rect 99840 3742 99892 3748
rect 99380 3392 99432 3398
rect 99380 3334 99432 3340
rect 99852 480 99880 3742
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100772 354 100800 11698
rect 102232 9036 102284 9042
rect 102232 8978 102284 8984
rect 102244 480 102272 8978
rect 104912 6914 104940 17206
rect 105556 11762 105584 38014
rect 106292 38010 106320 40063
rect 106660 40035 107100 40063
rect 106280 38004 106332 38010
rect 106280 37946 106332 37952
rect 106280 37392 106332 37398
rect 106280 37334 106332 37340
rect 106292 16574 106320 37334
rect 106660 26234 106688 40035
rect 106384 26206 106688 26234
rect 106384 25566 106412 26206
rect 106372 25560 106424 25566
rect 106372 25502 106424 25508
rect 106292 16546 106504 16574
rect 105544 11756 105596 11762
rect 105544 11698 105596 11704
rect 104912 6886 105768 6914
rect 104532 4888 104584 4894
rect 104532 4830 104584 4836
rect 103336 3868 103388 3874
rect 103336 3810 103388 3816
rect 103348 480 103376 3810
rect 104544 480 104572 4830
rect 105740 480 105768 6886
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 107672 11830 107700 40174
rect 108316 40066 108344 40174
rect 125612 40174 126284 40202
rect 107764 40035 107900 40063
rect 108316 40038 108680 40066
rect 109052 40035 109460 40063
rect 109788 40035 110240 40063
rect 110616 40035 111020 40063
rect 111800 40035 111840 40063
rect 107764 15978 107792 40035
rect 107752 15972 107804 15978
rect 107752 15914 107804 15920
rect 107660 11824 107712 11830
rect 107660 11766 107712 11772
rect 108120 4820 108172 4826
rect 108120 4762 108172 4768
rect 108132 480 108160 4762
rect 109052 3330 109080 40035
rect 109788 26234 109816 40035
rect 110420 37324 110472 37330
rect 110420 37266 110472 37272
rect 109144 26206 109816 26234
rect 109040 3324 109092 3330
rect 109040 3266 109092 3272
rect 109144 3262 109172 26206
rect 109316 7608 109368 7614
rect 109316 7550 109368 7556
rect 109132 3256 109184 3262
rect 109132 3198 109184 3204
rect 109328 480 109356 7550
rect 110432 6914 110460 37266
rect 110616 26234 110644 40035
rect 110524 26206 110644 26234
rect 110524 16574 110552 26206
rect 110524 16546 110644 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 110616 3738 110644 16546
rect 111616 13184 111668 13190
rect 111616 13126 111668 13132
rect 110604 3732 110656 3738
rect 110604 3674 110656 3680
rect 111628 480 111656 13126
rect 111812 3806 111840 40035
rect 112180 40035 112580 40063
rect 113284 40035 113360 40063
rect 114020 40035 114140 40063
rect 114572 40035 114900 40063
rect 115680 40035 115888 40063
rect 112180 26234 112208 40035
rect 113284 37398 113312 40035
rect 113272 37392 113324 37398
rect 113272 37334 113324 37340
rect 114020 37330 114048 40035
rect 114008 37324 114060 37330
rect 114008 37266 114060 37272
rect 111904 26206 112208 26234
rect 111904 3874 111932 26206
rect 112352 10396 112404 10402
rect 112352 10338 112404 10344
rect 111892 3868 111944 3874
rect 111892 3810 111944 3816
rect 111800 3800 111852 3806
rect 111800 3742 111852 3748
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 10338
rect 114572 2802 114600 40035
rect 115860 38010 115888 40035
rect 115952 40035 116460 40063
rect 116780 40035 117240 40063
rect 117700 40035 118040 40063
rect 118712 40035 118820 40063
rect 119172 40035 119600 40063
rect 120184 40035 120380 40063
rect 120736 40035 121160 40063
rect 121656 40035 121940 40063
rect 122300 40035 122720 40063
rect 123128 40035 123520 40063
rect 115848 38004 115900 38010
rect 115848 37946 115900 37952
rect 114744 14476 114796 14482
rect 114744 14418 114796 14424
rect 114480 2774 114600 2802
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 354 114090 480
rect 114480 354 114508 2774
rect 113978 326 114508 354
rect 114756 354 114784 14418
rect 115952 3126 115980 40035
rect 116780 38162 116808 40035
rect 116504 38134 116808 38162
rect 116504 26234 116532 38134
rect 116584 38004 116636 38010
rect 116584 37946 116636 37952
rect 116044 26206 116532 26234
rect 116044 3330 116072 26206
rect 116400 8968 116452 8974
rect 116400 8910 116452 8916
rect 116032 3324 116084 3330
rect 116032 3266 116084 3272
rect 115940 3120 115992 3126
rect 115940 3062 115992 3068
rect 116412 480 116440 8910
rect 116596 3534 116624 37946
rect 117700 26234 117728 40035
rect 117332 26206 117728 26234
rect 116584 3528 116636 3534
rect 116584 3470 116636 3476
rect 117332 3466 117360 26206
rect 118712 3602 118740 40035
rect 119172 26234 119200 40035
rect 118804 26206 119200 26234
rect 118804 16574 118832 26206
rect 118804 16546 119016 16574
rect 118792 6180 118844 6186
rect 118792 6122 118844 6128
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 117320 3460 117372 3466
rect 117320 3402 117372 3408
rect 117608 480 117636 3470
rect 118804 480 118832 6122
rect 118988 3670 119016 16546
rect 119896 11756 119948 11762
rect 119896 11698 119948 11704
rect 118976 3664 119028 3670
rect 118976 3606 119028 3612
rect 119908 480 119936 11698
rect 120184 3874 120212 40035
rect 120736 26234 120764 40035
rect 121656 37942 121684 40035
rect 121644 37936 121696 37942
rect 121644 37878 121696 37884
rect 121552 35216 121604 35222
rect 121552 35158 121604 35164
rect 120276 26206 120764 26234
rect 120172 3868 120224 3874
rect 120172 3810 120224 3816
rect 120276 3369 120304 26206
rect 121564 3482 121592 35158
rect 122300 26234 122328 40035
rect 122840 36644 122892 36650
rect 122840 36586 122892 36592
rect 121656 26206 122328 26234
rect 121656 3942 121684 26206
rect 121644 3936 121696 3942
rect 121644 3878 121696 3884
rect 121564 3454 122328 3482
rect 120262 3360 120318 3369
rect 120262 3295 120318 3304
rect 121092 3120 121144 3126
rect 121092 3062 121144 3068
rect 121104 480 121132 3062
rect 122300 480 122328 3454
rect 122852 490 122880 36586
rect 123128 26234 123156 40035
rect 124286 39794 124314 40049
rect 124784 40035 125080 40063
rect 124286 39766 124352 39794
rect 124220 38004 124272 38010
rect 124220 37946 124272 37952
rect 122944 26206 123156 26234
rect 122944 3262 122972 26206
rect 124232 3670 124260 37946
rect 124324 3738 124352 39766
rect 124784 38010 124812 40035
rect 124772 38004 124824 38010
rect 124772 37946 124824 37952
rect 124312 3732 124364 3738
rect 124312 3674 124364 3680
rect 124220 3664 124272 3670
rect 124220 3606 124272 3612
rect 125612 3466 125640 40174
rect 126256 40066 126284 40174
rect 136652 40174 137232 40202
rect 125704 40035 125860 40063
rect 126256 40038 126640 40066
rect 126992 40035 127400 40063
rect 128160 40035 128308 40063
rect 125600 3460 125652 3466
rect 125600 3402 125652 3408
rect 125704 3398 125732 40035
rect 125876 3936 125928 3942
rect 125876 3878 125928 3884
rect 125692 3392 125744 3398
rect 125692 3334 125744 3340
rect 124680 3324 124732 3330
rect 124680 3266 124732 3272
rect 122932 3256 122984 3262
rect 122932 3198 122984 3204
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 113978 -960 114090 326
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122852 462 123064 490
rect 124692 480 124720 3266
rect 125888 480 125916 3878
rect 126992 3602 127020 40035
rect 128280 38010 128308 40035
rect 128556 40035 128960 40063
rect 129740 40035 129780 40063
rect 130520 40035 130792 40063
rect 131300 40035 131620 40063
rect 132080 40035 132172 40063
rect 128268 38004 128320 38010
rect 128268 37946 128320 37952
rect 127072 35352 127124 35358
rect 127072 35294 127124 35300
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 127084 3482 127112 35294
rect 128556 26234 128584 40035
rect 129004 38004 129056 38010
rect 129004 37946 129056 37952
rect 128372 26206 128584 26234
rect 128372 8974 128400 26206
rect 129016 14550 129044 37946
rect 129752 21418 129780 40035
rect 130764 38078 130792 40035
rect 130752 38072 130804 38078
rect 130752 38014 130804 38020
rect 131592 37670 131620 40035
rect 132144 38010 132172 40035
rect 132512 40035 132860 40063
rect 133248 40035 133660 40063
rect 133984 40035 134440 40063
rect 134812 40035 135220 40063
rect 136000 40035 136312 40063
rect 132132 38004 132184 38010
rect 132132 37946 132184 37952
rect 131580 37664 131632 37670
rect 131580 37606 131632 37612
rect 129740 21412 129792 21418
rect 129740 21354 129792 21360
rect 129004 14544 129056 14550
rect 129004 14486 129056 14492
rect 129096 14476 129148 14482
rect 129096 14418 129148 14424
rect 128360 8968 128412 8974
rect 128360 8910 128412 8916
rect 129108 3534 129136 14418
rect 130568 11756 130620 11762
rect 130568 11698 130620 11704
rect 126992 3454 127112 3482
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 129096 3528 129148 3534
rect 129096 3470 129148 3476
rect 126992 480 127020 3454
rect 128188 480 128216 3470
rect 129372 3256 129424 3262
rect 129372 3198 129424 3204
rect 129384 480 129412 3198
rect 130580 480 130608 11698
rect 132512 10334 132540 40035
rect 133248 26234 133276 40035
rect 133788 37664 133840 37670
rect 133788 37606 133840 37612
rect 133800 36582 133828 37606
rect 133788 36576 133840 36582
rect 133788 36518 133840 36524
rect 133880 31340 133932 31346
rect 133880 31282 133932 31288
rect 132604 26206 133276 26234
rect 132604 13394 132632 26206
rect 132592 13388 132644 13394
rect 132592 13330 132644 13336
rect 132500 10328 132552 10334
rect 132500 10270 132552 10276
rect 131764 8084 131816 8090
rect 131764 8026 131816 8032
rect 131776 480 131804 8026
rect 132960 3732 133012 3738
rect 132960 3674 133012 3680
rect 132972 480 133000 3674
rect 123036 354 123064 462
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 31282
rect 133984 15978 134012 40035
rect 134812 26234 134840 40035
rect 136284 37942 136312 40035
rect 136272 37936 136324 37942
rect 136272 37878 136324 37884
rect 134076 26206 134840 26234
rect 134076 17270 134104 26206
rect 134064 17264 134116 17270
rect 134064 17206 134116 17212
rect 133972 15972 134024 15978
rect 133972 15914 134024 15920
rect 136652 5030 136680 40174
rect 137204 40066 137232 40174
rect 143644 40174 144224 40202
rect 136744 40035 136780 40063
rect 137204 40038 137560 40066
rect 138032 40035 138340 40063
rect 138676 40035 139120 40063
rect 139412 40035 139900 40063
rect 140332 40035 140680 40063
rect 141068 40035 141460 40063
rect 142220 40035 142292 40063
rect 136744 5098 136772 40035
rect 136824 17536 136876 17542
rect 136824 17478 136876 17484
rect 136836 16574 136864 17478
rect 136836 16546 137232 16574
rect 136732 5092 136784 5098
rect 136732 5034 136784 5040
rect 136640 5024 136692 5030
rect 136640 4966 136692 4972
rect 135260 3732 135312 3738
rect 135260 3674 135312 3680
rect 135272 480 135300 3674
rect 136456 3664 136508 3670
rect 136456 3606 136508 3612
rect 136468 480 136496 3606
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138032 4962 138060 40035
rect 138676 26234 138704 40035
rect 138124 26206 138704 26234
rect 138020 4956 138072 4962
rect 138020 4898 138072 4904
rect 138124 4894 138152 26206
rect 139412 18970 139440 40035
rect 140332 35894 140360 40035
rect 141068 35894 141096 40035
rect 141424 38072 141476 38078
rect 141424 38014 141476 38020
rect 142160 38072 142212 38078
rect 142160 38014 142212 38020
rect 139504 35866 140360 35894
rect 140792 35866 141096 35894
rect 139504 19990 139532 35866
rect 140044 27124 140096 27130
rect 140044 27066 140096 27072
rect 139492 19984 139544 19990
rect 139492 19926 139544 19932
rect 139400 18964 139452 18970
rect 139400 18906 139452 18912
rect 138848 13116 138900 13122
rect 138848 13058 138900 13064
rect 138112 4888 138164 4894
rect 138112 4830 138164 4836
rect 138860 480 138888 13058
rect 140056 3738 140084 27066
rect 140792 4826 140820 35866
rect 140872 34128 140924 34134
rect 140872 34070 140924 34076
rect 140884 16574 140912 34070
rect 140884 16546 141280 16574
rect 140780 4820 140832 4826
rect 140780 4762 140832 4768
rect 140044 3732 140096 3738
rect 140044 3674 140096 3680
rect 140044 3460 140096 3466
rect 140044 3402 140096 3408
rect 140056 480 140084 3402
rect 141252 480 141280 16546
rect 141436 7614 141464 38014
rect 141424 7608 141476 7614
rect 141424 7550 141476 7556
rect 142172 5302 142200 38014
rect 142264 5370 142292 40035
rect 142632 40035 143000 40063
rect 142632 38078 142660 40035
rect 142620 38072 142672 38078
rect 142620 38014 142672 38020
rect 143644 35894 143672 40174
rect 144196 40066 144224 40174
rect 157444 40174 158208 40202
rect 143766 39794 143794 40049
rect 144196 40038 144580 40066
rect 143552 35866 143672 35894
rect 143736 39766 143794 39794
rect 144932 40035 145360 40063
rect 145668 40035 146140 40063
rect 146496 40035 146920 40063
rect 143552 6526 143580 35866
rect 143632 31476 143684 31482
rect 143632 31418 143684 31424
rect 143644 16574 143672 31418
rect 143736 25838 143764 39766
rect 143724 25832 143776 25838
rect 143724 25774 143776 25780
rect 143644 16546 144776 16574
rect 143540 6520 143592 6526
rect 143540 6462 143592 6468
rect 142252 5364 142304 5370
rect 142252 5306 142304 5312
rect 142160 5296 142212 5302
rect 142160 5238 142212 5244
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 142436 3460 142488 3466
rect 142436 3402 142488 3408
rect 142448 480 142476 3402
rect 143552 480 143580 3470
rect 144748 480 144776 16546
rect 144932 6458 144960 40035
rect 145668 26234 145696 40035
rect 146496 26234 146524 40035
rect 146944 38004 146996 38010
rect 146944 37946 146996 37952
rect 145024 26206 145696 26234
rect 146312 26206 146524 26234
rect 144920 6452 144972 6458
rect 144920 6394 144972 6400
rect 145024 6390 145052 26206
rect 145012 6384 145064 6390
rect 145012 6326 145064 6332
rect 146312 6322 146340 26206
rect 146956 9042 146984 37946
rect 146944 9036 146996 9042
rect 146944 8978 146996 8984
rect 146300 6316 146352 6322
rect 146300 6258 146352 6264
rect 147692 6254 147720 40063
rect 148480 40035 148824 40063
rect 149280 40035 149560 40063
rect 148796 38010 148824 40035
rect 148784 38004 148836 38010
rect 148784 37946 148836 37952
rect 149532 37874 149560 40035
rect 149716 40035 150060 40063
rect 150452 40035 150840 40063
rect 151188 40035 151600 40063
rect 151832 40035 152380 40063
rect 152752 40035 153160 40063
rect 153580 40035 153940 40063
rect 149520 37868 149572 37874
rect 149520 37810 149572 37816
rect 149716 26234 149744 40035
rect 149072 26206 149744 26234
rect 149072 24546 149100 26206
rect 149060 24540 149112 24546
rect 149060 24482 149112 24488
rect 147864 15904 147916 15910
rect 147864 15846 147916 15852
rect 147680 6248 147732 6254
rect 147680 6190 147732 6196
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 145932 3528 145984 3534
rect 145932 3470 145984 3476
rect 145944 480 145972 3470
rect 147140 480 147168 3538
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 15846
rect 150452 6186 150480 40035
rect 151188 38026 151216 40035
rect 150544 37998 151216 38026
rect 150544 21554 150572 37998
rect 150624 37868 150676 37874
rect 150624 37810 150676 37816
rect 150636 32774 150664 37810
rect 150624 32768 150676 32774
rect 150624 32710 150676 32716
rect 151832 28422 151860 40035
rect 151820 28416 151872 28422
rect 151820 28358 151872 28364
rect 152752 26234 152780 40035
rect 153580 27062 153608 40035
rect 154726 39794 154754 40049
rect 155144 40035 155520 40063
rect 156280 40035 156552 40063
rect 154726 39766 154804 39794
rect 154672 38072 154724 38078
rect 154672 38014 154724 38020
rect 154580 36780 154632 36786
rect 154580 36722 154632 36728
rect 153568 27056 153620 27062
rect 153568 26998 153620 27004
rect 151924 26206 152780 26234
rect 151820 25968 151872 25974
rect 151820 25910 151872 25916
rect 150532 21548 150584 21554
rect 150532 21490 150584 21496
rect 150624 14544 150676 14550
rect 150624 14486 150676 14492
rect 150440 6180 150492 6186
rect 150440 6122 150492 6128
rect 149520 3596 149572 3602
rect 149520 3538 149572 3544
rect 149532 480 149560 3538
rect 150636 480 150664 14486
rect 151832 480 151860 25910
rect 151924 22914 151952 26206
rect 151912 22908 151964 22914
rect 151912 22850 151964 22856
rect 154212 8968 154264 8974
rect 154212 8910 154264 8916
rect 153016 3664 153068 3670
rect 153016 3606 153068 3612
rect 153028 480 153056 3606
rect 154224 480 154252 8910
rect 154592 6914 154620 36722
rect 154684 13258 154712 38014
rect 154776 29782 154804 39766
rect 155144 38078 155172 40035
rect 155132 38072 155184 38078
rect 155132 38014 155184 38020
rect 156524 36718 156552 40035
rect 156708 40035 157060 40063
rect 156512 36712 156564 36718
rect 156512 36654 156564 36660
rect 154764 29776 154816 29782
rect 154764 29718 154816 29724
rect 156708 26234 156736 40035
rect 155972 26206 156736 26234
rect 155972 14550 156000 26206
rect 157340 21412 157392 21418
rect 157340 21354 157392 21360
rect 157352 16574 157380 21354
rect 157444 18766 157472 40174
rect 158180 40066 158208 40174
rect 160112 40174 160600 40202
rect 157536 40035 157840 40063
rect 158180 40038 158620 40066
rect 159008 40035 159400 40063
rect 157536 20126 157564 40035
rect 158720 29980 158772 29986
rect 158720 29922 158772 29928
rect 157524 20120 157576 20126
rect 157524 20062 157576 20068
rect 157432 18760 157484 18766
rect 157432 18702 157484 18708
rect 158732 16574 158760 29922
rect 159008 26234 159036 40035
rect 158824 26206 159036 26234
rect 158824 25702 158852 26206
rect 158812 25696 158864 25702
rect 158812 25638 158864 25644
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 155960 14544 156012 14550
rect 155960 14486 156012 14492
rect 154672 13252 154724 13258
rect 154672 13194 154724 13200
rect 154592 6886 155448 6914
rect 155420 480 155448 6886
rect 156604 3732 156656 3738
rect 156604 3674 156656 3680
rect 156616 480 156644 3674
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 7750 160140 40174
rect 160572 40066 160600 40174
rect 161584 40174 162164 40202
rect 160200 40035 160232 40063
rect 160572 40038 160980 40066
rect 160204 32638 160232 40035
rect 161480 34196 161532 34202
rect 161480 34138 161532 34144
rect 160192 32632 160244 32638
rect 160192 32574 160244 32580
rect 160100 7744 160152 7750
rect 160100 7686 160152 7692
rect 161296 7608 161348 7614
rect 161296 7550 161348 7556
rect 160100 3800 160152 3806
rect 160100 3742 160152 3748
rect 160112 480 160140 3742
rect 161308 480 161336 7550
rect 161492 6914 161520 34138
rect 161584 7614 161612 40174
rect 162136 40066 162164 40174
rect 172532 40174 173112 40202
rect 161676 40035 161760 40063
rect 162136 40038 162540 40066
rect 163320 40035 163636 40063
rect 161676 7682 161704 40035
rect 163608 38214 163636 40035
rect 163700 40035 164100 40063
rect 164436 40035 164880 40063
rect 165660 40035 165752 40063
rect 163596 38208 163648 38214
rect 163596 38150 163648 38156
rect 163700 33998 163728 40035
rect 164240 36576 164292 36582
rect 164240 36518 164292 36524
rect 163688 33992 163740 33998
rect 163688 33934 163740 33940
rect 164252 16574 164280 36518
rect 164436 26234 164464 40035
rect 165620 38072 165672 38078
rect 165620 38014 165672 38020
rect 164344 26206 164464 26234
rect 164344 21622 164372 26206
rect 165632 22982 165660 38014
rect 165724 28558 165752 40035
rect 166184 40035 166440 40063
rect 167220 40035 167500 40063
rect 166184 38078 166212 40035
rect 166172 38072 166224 38078
rect 166172 38014 166224 38020
rect 167472 36854 167500 40035
rect 167564 40035 168000 40063
rect 168392 40035 168780 40063
rect 169560 40035 169708 40063
rect 167460 36848 167512 36854
rect 167460 36790 167512 36796
rect 167000 35488 167052 35494
rect 167000 35430 167052 35436
rect 165712 28552 165764 28558
rect 165712 28494 165764 28500
rect 165620 22976 165672 22982
rect 165620 22918 165672 22924
rect 164332 21616 164384 21622
rect 164332 21558 164384 21564
rect 167012 16574 167040 35430
rect 167564 27198 167592 40035
rect 168392 29850 168420 40035
rect 169680 38146 169708 40035
rect 169956 40035 170340 40063
rect 171120 40035 171364 40063
rect 169668 38140 169720 38146
rect 169668 38082 169720 38088
rect 168380 29844 168432 29850
rect 168380 29786 168432 29792
rect 167552 27192 167604 27198
rect 167552 27134 167604 27140
rect 169956 26234 169984 40035
rect 171336 38214 171364 40035
rect 171428 40035 171900 40063
rect 170404 38208 170456 38214
rect 170404 38150 170456 38156
rect 171324 38208 171376 38214
rect 171324 38150 171376 38156
rect 169772 26206 169984 26234
rect 169772 17474 169800 26206
rect 170416 24274 170444 38150
rect 171428 35426 171456 40035
rect 171416 35420 171468 35426
rect 171416 35362 171468 35368
rect 170404 24268 170456 24274
rect 170404 24210 170456 24216
rect 169760 17468 169812 17474
rect 169760 17410 169812 17416
rect 164252 16546 164464 16574
rect 167012 16546 167224 16574
rect 163688 13184 163740 13190
rect 163688 13126 163740 13132
rect 161664 7676 161716 7682
rect 161664 7618 161716 7624
rect 161572 7608 161624 7614
rect 161572 7550 161624 7556
rect 161492 6886 162072 6914
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 6886
rect 163700 480 163728 13126
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166080 13320 166132 13326
rect 166080 13262 166132 13268
rect 166092 480 166120 13262
rect 167196 480 167224 16546
rect 170312 14816 170364 14822
rect 170312 14758 170364 14764
rect 168380 11824 168432 11830
rect 168380 11766 168432 11772
rect 168392 3874 168420 11766
rect 168472 9036 168524 9042
rect 168472 8978 168524 8984
rect 168380 3868 168432 3874
rect 168380 3810 168432 3816
rect 168484 3482 168512 8978
rect 169576 3868 169628 3874
rect 169576 3810 169628 3816
rect 168392 3454 168512 3482
rect 168392 480 168420 3454
rect 169588 480 169616 3810
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 14758
rect 171968 10328 172020 10334
rect 171968 10270 172020 10276
rect 171980 480 172008 10270
rect 172532 9586 172560 40174
rect 173084 40066 173112 40174
rect 173912 40174 174584 40202
rect 172666 39794 172694 40049
rect 173084 40038 173460 40066
rect 172624 39766 172694 39794
rect 172624 18834 172652 39766
rect 172704 38208 172756 38214
rect 172704 38150 172756 38156
rect 172716 31278 172744 38150
rect 172704 31272 172756 31278
rect 172704 31214 172756 31220
rect 172612 18828 172664 18834
rect 172612 18770 172664 18776
rect 172704 11892 172756 11898
rect 172704 11834 172756 11840
rect 172520 9580 172572 9586
rect 172520 9522 172572 9528
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 11834
rect 173912 9450 173940 40174
rect 174556 40066 174584 40174
rect 190472 40174 191052 40202
rect 174004 40035 174240 40063
rect 174556 40038 175020 40066
rect 175292 40035 175800 40063
rect 176212 40035 176580 40063
rect 176948 40035 177360 40063
rect 178052 40035 178140 40063
rect 178512 40035 178920 40063
rect 179432 40035 179700 40063
rect 180076 40035 180500 40063
rect 181280 40035 181576 40063
rect 174004 9518 174032 40035
rect 174084 18896 174136 18902
rect 174084 18838 174136 18844
rect 173992 9512 174044 9518
rect 173992 9454 174044 9460
rect 173900 9444 173952 9450
rect 173900 9386 173952 9392
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 174096 354 174124 18838
rect 175292 9382 175320 40035
rect 176212 26234 176240 40035
rect 176948 35894 176976 40035
rect 177304 37936 177356 37942
rect 177304 37878 177356 37884
rect 175384 26206 176240 26234
rect 176672 35866 176976 35894
rect 175280 9376 175332 9382
rect 175280 9318 175332 9324
rect 175384 9314 175412 26206
rect 175464 13388 175516 13394
rect 175464 13330 175516 13336
rect 175372 9308 175424 9314
rect 175372 9250 175424 9256
rect 175476 480 175504 13330
rect 176672 9246 176700 35866
rect 176752 28484 176804 28490
rect 176752 28426 176804 28432
rect 176660 9240 176712 9246
rect 176660 9182 176712 9188
rect 176764 3874 176792 28426
rect 176844 11960 176896 11966
rect 176844 11902 176896 11908
rect 176752 3868 176804 3874
rect 176752 3810 176804 3816
rect 176856 3482 176884 11902
rect 177316 10334 177344 37878
rect 177304 10328 177356 10334
rect 177304 10270 177356 10276
rect 178052 9178 178080 40035
rect 178512 26234 178540 40035
rect 178144 26206 178540 26234
rect 178040 9172 178092 9178
rect 178040 9114 178092 9120
rect 178144 9110 178172 26206
rect 178592 15972 178644 15978
rect 178592 15914 178644 15920
rect 178132 9104 178184 9110
rect 178132 9046 178184 9052
rect 177856 3868 177908 3874
rect 177856 3810 177908 3816
rect 176672 3454 176884 3482
rect 176672 480 176700 3454
rect 177868 480 177896 3810
rect 174238 354 174350 480
rect 174096 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 15914
rect 179432 9042 179460 40035
rect 180076 26234 180104 40035
rect 181548 38214 181576 40035
rect 181640 40035 182060 40063
rect 182468 40035 182840 40063
rect 181536 38208 181588 38214
rect 181536 38150 181588 38156
rect 181640 32570 181668 40035
rect 181628 32564 181680 32570
rect 181628 32506 181680 32512
rect 182468 26234 182496 40035
rect 183606 39794 183634 40049
rect 179524 26206 180104 26234
rect 182192 26206 182496 26234
rect 183572 39766 183634 39794
rect 183940 40035 184400 40063
rect 185160 40035 185440 40063
rect 185960 40035 186268 40063
rect 186740 40035 187004 40063
rect 179420 9036 179472 9042
rect 179420 8978 179472 8984
rect 179524 8974 179552 26206
rect 182192 24342 182220 26206
rect 182180 24336 182232 24342
rect 182180 24278 182232 24284
rect 183572 21486 183600 39766
rect 183940 28354 183968 40035
rect 185412 38282 185440 40035
rect 185400 38276 185452 38282
rect 185400 38218 185452 38224
rect 186240 36582 186268 40035
rect 186976 37942 187004 40035
rect 187068 40035 187520 40063
rect 187896 40035 188300 40063
rect 189060 40035 189212 40063
rect 186964 37936 187016 37942
rect 186964 37878 187016 37884
rect 186228 36576 186280 36582
rect 186228 36518 186280 36524
rect 183928 28348 183980 28354
rect 183928 28290 183980 28296
rect 187068 26994 187096 40035
rect 187056 26988 187108 26994
rect 187056 26930 187108 26936
rect 187896 26234 187924 40035
rect 188344 38276 188396 38282
rect 188344 38218 188396 38224
rect 187712 26206 187924 26234
rect 184940 24404 184992 24410
rect 184940 24346 184992 24352
rect 183560 21480 183612 21486
rect 183560 21422 183612 21428
rect 182180 17264 182232 17270
rect 182180 17206 182232 17212
rect 180984 15972 181036 15978
rect 180984 15914 181036 15920
rect 180248 12028 180300 12034
rect 180248 11970 180300 11976
rect 179512 8968 179564 8974
rect 179512 8910 179564 8916
rect 180260 480 180288 11970
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 15914
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 17206
rect 183744 12096 183796 12102
rect 183744 12038 183796 12044
rect 183756 480 183784 12038
rect 184952 480 184980 24346
rect 186872 12164 186924 12170
rect 186872 12106 186924 12112
rect 186136 10328 186188 10334
rect 186136 10270 186188 10276
rect 186148 480 186176 10270
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 12106
rect 187712 10674 187740 26206
rect 188356 22846 188384 38218
rect 189184 37670 189212 40035
rect 189460 40035 189840 40063
rect 189172 37664 189224 37670
rect 189172 37606 189224 37612
rect 189460 26234 189488 40035
rect 189092 26206 189488 26234
rect 188344 22840 188396 22846
rect 188344 22782 188396 22788
rect 189092 20058 189120 26206
rect 189080 20052 189132 20058
rect 189080 19994 189132 20000
rect 188528 16108 188580 16114
rect 188528 16050 188580 16056
rect 187700 10668 187752 10674
rect 187700 10610 187752 10616
rect 188540 480 188568 16050
rect 190472 10538 190500 40174
rect 191024 40066 191052 40174
rect 191852 40174 192616 40202
rect 190606 39794 190634 40049
rect 191024 40038 191420 40066
rect 190564 39766 190634 39794
rect 190564 10606 190592 39766
rect 190644 37664 190696 37670
rect 190644 37606 190696 37612
rect 190656 29714 190684 37606
rect 190644 29708 190696 29714
rect 190644 29650 190696 29656
rect 190644 12232 190696 12238
rect 190644 12174 190696 12180
rect 190552 10600 190604 10606
rect 190552 10542 190604 10548
rect 190460 10532 190512 10538
rect 190460 10474 190512 10480
rect 189724 5092 189776 5098
rect 189724 5034 189776 5040
rect 189736 480 189764 5034
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190656 354 190684 12174
rect 191852 10402 191880 40174
rect 192588 40066 192616 40174
rect 195992 40174 196480 40202
rect 191944 40035 192200 40063
rect 192588 40038 192980 40066
rect 193760 40035 194088 40063
rect 191944 10470 191972 40035
rect 194060 38486 194088 40035
rect 194152 40035 194540 40063
rect 194980 40035 195320 40063
rect 194048 38480 194100 38486
rect 194048 38422 194100 38428
rect 194152 26234 194180 40035
rect 194980 26234 195008 40035
rect 195244 38480 195296 38486
rect 195244 38422 195296 38428
rect 193232 26206 194180 26234
rect 194612 26206 195008 26234
rect 193232 25634 193260 26206
rect 193220 25628 193272 25634
rect 193220 25570 193272 25576
rect 192024 16176 192076 16182
rect 192024 16118 192076 16124
rect 191932 10464 191984 10470
rect 191932 10406 191984 10412
rect 191840 10396 191892 10402
rect 191840 10338 191892 10344
rect 192036 480 192064 16118
rect 193220 14612 193272 14618
rect 193220 14554 193272 14560
rect 193232 3398 193260 14554
rect 194612 10334 194640 26206
rect 194692 23044 194744 23050
rect 194692 22986 194744 22992
rect 194704 16574 194732 22986
rect 195256 18698 195284 38422
rect 195244 18692 195296 18698
rect 195244 18634 195296 18640
rect 195992 17406 196020 40174
rect 196452 40066 196480 40174
rect 197372 40174 198136 40202
rect 196084 40035 196120 40063
rect 196452 40038 196900 40066
rect 196084 33930 196112 40035
rect 196072 33924 196124 33930
rect 196072 33866 196124 33872
rect 197372 24206 197400 40174
rect 198108 40066 198136 40174
rect 208412 40174 208992 40202
rect 197464 40035 197680 40063
rect 198108 40038 198460 40066
rect 199220 40035 199516 40063
rect 197464 32502 197492 40035
rect 199488 38078 199516 40035
rect 199580 40035 200000 40063
rect 200316 40035 200780 40063
rect 199476 38072 199528 38078
rect 199476 38014 199528 38020
rect 197452 32496 197504 32502
rect 197452 32438 197504 32444
rect 199580 31210 199608 40035
rect 199568 31204 199620 31210
rect 199568 31146 199620 31152
rect 200316 26234 200344 40035
rect 201546 39794 201574 40049
rect 201512 39766 201574 39794
rect 201972 40035 202340 40063
rect 203120 40035 203472 40063
rect 203900 40035 204208 40063
rect 200764 38140 200816 38146
rect 200764 38082 200816 38088
rect 200132 26206 200344 26234
rect 197360 24200 197412 24206
rect 197360 24142 197412 24148
rect 195980 17400 196032 17406
rect 195980 17342 196032 17348
rect 200132 17338 200160 26206
rect 200776 20194 200804 38082
rect 201512 35290 201540 39766
rect 201500 35284 201552 35290
rect 201500 35226 201552 35232
rect 201972 26234 202000 40035
rect 203444 38282 203472 40035
rect 203432 38276 203484 38282
rect 203432 38218 203484 38224
rect 204180 37874 204208 40035
rect 204364 40035 204680 40063
rect 205100 40035 205460 40063
rect 205836 40035 206240 40063
rect 207040 40035 207336 40063
rect 204168 37868 204220 37874
rect 204168 37810 204220 37816
rect 204260 35556 204312 35562
rect 204260 35498 204312 35504
rect 201604 26206 202000 26234
rect 201500 25900 201552 25906
rect 201500 25842 201552 25848
rect 200764 20188 200816 20194
rect 200764 20130 200816 20136
rect 200120 17332 200172 17338
rect 200120 17274 200172 17280
rect 194704 16546 195192 16574
rect 194600 10328 194652 10334
rect 194600 10270 194652 10276
rect 193312 5024 193364 5030
rect 193312 4966 193364 4972
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 193324 2530 193352 4966
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 193232 2502 193352 2530
rect 193232 480 193260 2502
rect 194428 480 194456 3334
rect 190798 354 190910 480
rect 190656 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 198740 16312 198792 16318
rect 198740 16254 198792 16260
rect 197912 12300 197964 12306
rect 197912 12242 197964 12248
rect 196808 4956 196860 4962
rect 196808 4898 196860 4904
rect 196820 480 196848 4898
rect 197924 480 197952 12242
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 16254
rect 201512 11694 201540 25842
rect 201604 18630 201632 26206
rect 202880 18964 202932 18970
rect 202880 18906 202932 18912
rect 201592 18624 201644 18630
rect 201592 18566 201644 18572
rect 202892 16574 202920 18906
rect 204272 16574 204300 35498
rect 204364 21418 204392 40035
rect 205100 29646 205128 40035
rect 205640 29912 205692 29918
rect 205640 29854 205692 29860
rect 205088 29640 205140 29646
rect 205088 29582 205140 29588
rect 204352 21412 204404 21418
rect 204352 21354 204404 21360
rect 205652 16574 205680 29854
rect 205836 26234 205864 40035
rect 207308 38418 207336 40035
rect 207400 40035 207820 40063
rect 207296 38412 207348 38418
rect 207296 38354 207348 38360
rect 206928 37868 206980 37874
rect 206928 37810 206980 37816
rect 206940 31142 206968 37810
rect 206928 31136 206980 31142
rect 206928 31078 206980 31084
rect 207400 26926 207428 40035
rect 207388 26920 207440 26926
rect 207388 26862 207440 26868
rect 205744 26206 205864 26234
rect 205744 22778 205772 26206
rect 205732 22772 205784 22778
rect 205732 22714 205784 22720
rect 207020 19984 207072 19990
rect 207020 19926 207072 19932
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 201592 13388 201644 13394
rect 201592 13330 201644 13336
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 13330
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 200304 4888 200356 4894
rect 200304 4830 200356 4836
rect 200316 480 200344 4830
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 19926
rect 208412 5166 208440 40174
rect 208964 40066 208992 40174
rect 209884 40174 210556 40202
rect 208504 40035 208600 40063
rect 208964 40038 209380 40066
rect 208504 5234 208532 40035
rect 209044 38412 209096 38418
rect 209044 38354 209096 38360
rect 209056 28286 209084 38354
rect 209884 35894 209912 40174
rect 210528 40066 210556 40174
rect 234724 40174 235488 40202
rect 209792 35866 209912 35894
rect 209976 40035 210160 40063
rect 210528 40038 210940 40066
rect 211356 40035 211740 40063
rect 212520 40035 212764 40063
rect 209044 28280 209096 28286
rect 209044 28222 209096 28228
rect 208584 7812 208636 7818
rect 208584 7754 208636 7760
rect 208492 5228 208544 5234
rect 208492 5170 208544 5176
rect 208400 5160 208452 5166
rect 208400 5102 208452 5108
rect 208596 480 208624 7754
rect 209792 5098 209820 35866
rect 209872 34060 209924 34066
rect 209872 34002 209924 34008
rect 209780 5092 209832 5098
rect 209780 5034 209832 5040
rect 209884 3482 209912 34002
rect 209976 24138 210004 40035
rect 211356 26234 211384 40035
rect 212540 39568 212592 39574
rect 212540 39510 212592 39516
rect 211172 26206 211384 26234
rect 209964 24132 210016 24138
rect 209964 24074 210016 24080
rect 211172 5030 211200 26206
rect 211712 14680 211764 14686
rect 211712 14622 211764 14628
rect 211160 5024 211212 5030
rect 211160 4966 211212 4972
rect 210976 4820 211028 4826
rect 210976 4762 211028 4768
rect 209792 3454 209912 3482
rect 209792 480 209820 3454
rect 210988 480 211016 4762
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 14622
rect 212552 4894 212580 39510
rect 212736 26234 212764 40035
rect 212920 40035 213280 40063
rect 213932 40035 214040 40063
rect 214392 40035 214820 40063
rect 215600 40035 215892 40063
rect 212920 39574 212948 40035
rect 212908 39568 212960 39574
rect 212908 39510 212960 39516
rect 212644 26206 212764 26234
rect 212644 4962 212672 26206
rect 212724 17604 212776 17610
rect 212724 17546 212776 17552
rect 212736 16574 212764 17546
rect 212736 16546 213408 16574
rect 212632 4956 212684 4962
rect 212632 4898 212684 4904
rect 212540 4888 212592 4894
rect 212540 4830 212592 4836
rect 213380 480 213408 16546
rect 213932 4758 213960 40035
rect 214392 26234 214420 40035
rect 215864 38146 215892 40035
rect 215956 40035 216380 40063
rect 216784 40035 217180 40063
rect 217888 40038 217960 40066
rect 215852 38140 215904 38146
rect 215852 38082 215904 38088
rect 215956 26234 215984 40035
rect 216784 32434 216812 40035
rect 217324 38004 217376 38010
rect 217324 37946 217376 37952
rect 216772 32428 216824 32434
rect 216772 32370 216824 32376
rect 216680 31408 216732 31414
rect 216680 31350 216732 31356
rect 214024 26206 214420 26234
rect 215312 26206 215984 26234
rect 214024 25566 214052 26206
rect 214012 25560 214064 25566
rect 214012 25502 214064 25508
rect 215312 19990 215340 26206
rect 215300 19984 215352 19990
rect 215300 19926 215352 19932
rect 216692 16574 216720 31350
rect 216692 16546 216904 16574
rect 215300 13456 215352 13462
rect 215300 13398 215352 13404
rect 214472 5364 214524 5370
rect 214472 5306 214524 5312
rect 213920 4752 213972 4758
rect 213920 4694 213972 4700
rect 214484 480 214512 5306
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 13398
rect 216876 480 216904 16546
rect 217336 13530 217364 37946
rect 217888 36650 217916 40038
rect 218740 40035 218836 40063
rect 218704 38208 218756 38214
rect 218704 38150 218756 38156
rect 217876 36644 217928 36650
rect 217876 36586 217928 36592
rect 218716 25770 218744 38150
rect 218808 38010 218836 40035
rect 219506 39794 219534 40049
rect 220004 40035 220300 40063
rect 220832 40035 221080 40063
rect 221860 40035 222148 40063
rect 219506 39766 219572 39794
rect 218796 38004 218848 38010
rect 218796 37946 218848 37952
rect 219440 37868 219492 37874
rect 219440 37810 219492 37816
rect 218704 25764 218756 25770
rect 218704 25706 218756 25712
rect 219452 17270 219480 37810
rect 219544 35222 219572 39766
rect 220004 37874 220032 40035
rect 219992 37868 220044 37874
rect 219992 37810 220044 37816
rect 219532 35216 219584 35222
rect 219532 35158 219584 35164
rect 220832 33794 220860 40035
rect 222120 37874 222148 40035
rect 222212 40035 222660 40063
rect 223040 40035 223440 40063
rect 223868 40035 224220 40063
rect 222108 37868 222160 37874
rect 222108 37810 222160 37816
rect 222212 35358 222240 40035
rect 223040 38842 223068 40035
rect 222580 38814 223068 38842
rect 222580 35894 222608 38814
rect 222660 37868 222712 37874
rect 222660 37810 222712 37816
rect 222304 35866 222608 35894
rect 222200 35352 222252 35358
rect 222200 35294 222252 35300
rect 220820 33788 220872 33794
rect 220820 33730 220872 33736
rect 220820 25832 220872 25838
rect 220820 25774 220872 25780
rect 219532 21752 219584 21758
rect 219532 21694 219584 21700
rect 219440 17264 219492 17270
rect 219440 17206 219492 17212
rect 219544 16574 219572 21694
rect 220832 16574 220860 25774
rect 219544 16546 220032 16574
rect 220832 16546 221136 16574
rect 218060 14748 218112 14754
rect 218060 14690 218112 14696
rect 217324 13524 217376 13530
rect 217324 13466 217376 13472
rect 218072 7546 218100 14690
rect 218060 7540 218112 7546
rect 218060 7482 218112 7488
rect 219256 7540 219308 7546
rect 219256 7482 219308 7488
rect 218152 5296 218204 5302
rect 218152 5238 218204 5244
rect 218164 2666 218192 5238
rect 218072 2638 218192 2666
rect 218072 480 218100 2638
rect 219268 480 219296 7482
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222304 11762 222332 35866
rect 222384 35624 222436 35630
rect 222384 35566 222436 35572
rect 222396 16574 222424 35566
rect 222672 31074 222700 37810
rect 223580 36916 223632 36922
rect 223580 36858 223632 36864
rect 222660 31068 222712 31074
rect 222660 31010 222712 31016
rect 222396 16546 222792 16574
rect 222292 11756 222344 11762
rect 222292 11698 222344 11704
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 36858
rect 223868 31346 223896 40035
rect 224132 38276 224184 38282
rect 224132 38218 224184 38224
rect 224144 33862 224172 38218
rect 224972 37874 225000 40063
rect 225340 40035 225760 40063
rect 226352 40035 226540 40063
rect 226996 40035 227340 40063
rect 227824 40035 228100 40063
rect 228560 40035 228880 40063
rect 229204 40035 229660 40063
rect 230032 40035 230440 40063
rect 230860 40035 231220 40063
rect 231872 40035 232000 40063
rect 232332 40035 232800 40063
rect 233252 40035 233580 40063
rect 233988 40035 234360 40063
rect 224224 37868 224276 37874
rect 224224 37810 224276 37816
rect 224960 37868 225012 37874
rect 224960 37810 225012 37816
rect 224132 33856 224184 33862
rect 224132 33798 224184 33804
rect 223856 31340 223908 31346
rect 223856 31282 223908 31288
rect 224236 17542 224264 37810
rect 225340 34134 225368 40035
rect 225328 34128 225380 34134
rect 225328 34070 225380 34076
rect 226352 31482 226380 40035
rect 226996 38570 227024 40035
rect 226536 38542 227024 38570
rect 226340 31476 226392 31482
rect 226340 31418 226392 31424
rect 226536 26234 226564 38542
rect 226616 38208 226668 38214
rect 226616 38150 226668 38156
rect 226444 26206 226564 26234
rect 224224 17536 224276 17542
rect 224224 17478 224276 17484
rect 226444 15910 226472 26206
rect 226432 15904 226484 15910
rect 226432 15846 226484 15852
rect 226628 6914 226656 38150
rect 227824 25974 227852 40035
rect 228560 36786 228588 40035
rect 229204 39794 229232 40035
rect 229112 39766 229232 39794
rect 228548 36780 228600 36786
rect 228548 36722 228600 36728
rect 229112 29986 229140 39766
rect 230032 34202 230060 40035
rect 230020 34196 230072 34202
rect 230020 34138 230072 34144
rect 229100 29980 229152 29986
rect 229100 29922 229152 29928
rect 230860 26234 230888 40035
rect 230492 26206 230888 26234
rect 227812 25968 227864 25974
rect 227812 25910 227864 25916
rect 227536 16380 227588 16386
rect 227536 16322 227588 16328
rect 226352 6886 226656 6914
rect 225144 6520 225196 6526
rect 225144 6462 225196 6468
rect 225156 480 225184 6462
rect 226352 480 226380 6886
rect 227548 480 227576 16322
rect 230492 13326 230520 26206
rect 231032 14884 231084 14890
rect 231032 14826 231084 14832
rect 230480 13320 230532 13326
rect 230480 13262 230532 13268
rect 228732 6452 228784 6458
rect 228732 6394 228784 6400
rect 229836 6452 229888 6458
rect 229836 6394 229888 6400
rect 228744 480 228772 6394
rect 229848 480 229876 6394
rect 231044 480 231072 14826
rect 231872 11830 231900 40035
rect 232332 26234 232360 40035
rect 231964 26206 232360 26234
rect 231964 11898 231992 26206
rect 233252 11966 233280 40035
rect 233988 26234 234016 40035
rect 234620 32700 234672 32706
rect 234620 32642 234672 32648
rect 233344 26206 234016 26234
rect 233344 12034 233372 26206
rect 233332 12028 233384 12034
rect 233332 11970 233384 11976
rect 233240 11960 233292 11966
rect 233240 11902 233292 11908
rect 231952 11892 232004 11898
rect 231952 11834 232004 11840
rect 231860 11824 231912 11830
rect 231860 11766 231912 11772
rect 233424 11756 233476 11762
rect 233424 11698 233476 11704
rect 232228 6384 232280 6390
rect 232228 6326 232280 6332
rect 232240 480 232268 6326
rect 233436 480 233464 11698
rect 234632 480 234660 32642
rect 234724 12170 234752 40174
rect 235460 40066 235488 40174
rect 237392 40174 237880 40202
rect 234816 40035 235140 40063
rect 235460 40038 235920 40066
rect 236288 40035 236700 40063
rect 234712 12164 234764 12170
rect 234712 12106 234764 12112
rect 234816 12102 234844 40035
rect 236288 26234 236316 40035
rect 236012 26206 236316 26234
rect 236012 12238 236040 26206
rect 237392 12306 237420 40174
rect 237852 40066 237880 40174
rect 255332 40174 255820 40202
rect 237480 40035 237512 40063
rect 237852 40038 238260 40066
rect 237484 14618 237512 40035
rect 238772 40035 239040 40063
rect 239416 40035 239820 40063
rect 240152 40035 240600 40063
rect 240980 40035 241380 40063
rect 241716 40035 242160 40063
rect 237564 20256 237616 20262
rect 237564 20198 237616 20204
rect 237576 16574 237604 20198
rect 237576 16546 237696 16574
rect 237472 14612 237524 14618
rect 237472 14554 237524 14560
rect 237380 12300 237432 12306
rect 237380 12242 237432 12248
rect 236000 12232 236052 12238
rect 236000 12174 236052 12180
rect 234804 12096 234856 12102
rect 234804 12038 234856 12044
rect 236552 11824 236604 11830
rect 236552 11766 236604 11772
rect 235816 6316 235868 6322
rect 235816 6258 235868 6264
rect 235828 480 235856 6258
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 11766
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 238772 13394 238800 40035
rect 239416 35562 239444 40035
rect 239404 35556 239456 35562
rect 239404 35498 239456 35504
rect 238760 13388 238812 13394
rect 238760 13330 238812 13336
rect 240152 7818 240180 40035
rect 240980 26234 241008 40035
rect 241716 26234 241744 40035
rect 242912 37874 242940 40063
rect 243372 40035 243720 40063
rect 244292 40035 244500 40063
rect 244844 40035 245280 40063
rect 245764 40035 246060 40063
rect 246500 40035 246840 40063
rect 247236 40035 247620 40063
rect 248420 40035 248552 40063
rect 242164 37868 242216 37874
rect 242164 37810 242216 37816
rect 242900 37868 242952 37874
rect 242900 37810 242952 37816
rect 240244 26206 241008 26234
rect 241532 26206 241744 26234
rect 240244 14686 240272 26206
rect 240232 14680 240284 14686
rect 240232 14622 240284 14628
rect 241532 13462 241560 26206
rect 241612 24472 241664 24478
rect 241612 24414 241664 24420
rect 241624 16574 241652 24414
rect 241624 16546 241744 16574
rect 241520 13456 241572 13462
rect 241520 13398 241572 13404
rect 240232 11416 240284 11422
rect 240232 11358 240284 11364
rect 240140 7812 240192 7818
rect 240140 7754 240192 7760
rect 239312 6248 239364 6254
rect 239312 6190 239364 6196
rect 239324 480 239352 6190
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240244 354 240272 11358
rect 241716 480 241744 16546
rect 242176 14754 242204 37810
rect 243372 35630 243400 40035
rect 244292 38214 244320 40035
rect 244280 38208 244332 38214
rect 244280 38150 244332 38156
rect 243360 35624 243412 35630
rect 243360 35566 243412 35572
rect 244372 29980 244424 29986
rect 244372 29922 244424 29928
rect 242164 14748 242216 14754
rect 242164 14690 242216 14696
rect 242900 13524 242952 13530
rect 242900 13466 242952 13472
rect 242912 480 242940 13466
rect 244096 5636 244148 5642
rect 244096 5578 244148 5584
rect 244108 480 244136 5578
rect 244384 3482 244412 29922
rect 244844 26234 244872 40035
rect 245764 37874 245792 40035
rect 244924 37868 244976 37874
rect 244924 37810 244976 37816
rect 245752 37868 245804 37874
rect 245752 37810 245804 37816
rect 244476 26206 244872 26234
rect 244476 6458 244504 26206
rect 244936 11762 244964 37810
rect 245660 32768 245712 32774
rect 245660 32710 245712 32716
rect 244924 11756 244976 11762
rect 244924 11698 244976 11704
rect 245672 6914 245700 32710
rect 246500 26234 246528 40035
rect 247236 26234 247264 40035
rect 248420 37868 248472 37874
rect 248420 37810 248472 37816
rect 245764 26206 246528 26234
rect 247052 26206 247264 26234
rect 245764 11830 245792 26206
rect 245752 11824 245804 11830
rect 245752 11766 245804 11772
rect 247052 11422 247080 26206
rect 247040 11416 247092 11422
rect 247040 11358 247092 11364
rect 245672 6886 245976 6914
rect 244464 6452 244516 6458
rect 244464 6394 244516 6400
rect 244384 3454 245240 3482
rect 245212 480 245240 3454
rect 240478 354 240590 480
rect 240244 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 6886
rect 248432 5574 248460 37810
rect 248524 5642 248552 40035
rect 248892 40035 249200 40063
rect 249812 40035 249960 40063
rect 250364 40035 250740 40063
rect 251284 40035 251520 40063
rect 251836 40035 252300 40063
rect 252664 40035 253080 40063
rect 253584 40035 253880 40063
rect 254228 40035 254660 40063
rect 248892 37874 248920 40035
rect 248880 37868 248932 37874
rect 248880 37810 248932 37816
rect 248604 25968 248656 25974
rect 248604 25910 248656 25916
rect 248512 5636 248564 5642
rect 248512 5578 248564 5584
rect 247592 5568 247644 5574
rect 247592 5510 247644 5516
rect 248420 5568 248472 5574
rect 248420 5510 248472 5516
rect 247604 480 247632 5510
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248616 354 248644 25910
rect 249812 11898 249840 40035
rect 250364 26234 250392 40035
rect 251180 35624 251232 35630
rect 251180 35566 251232 35572
rect 249904 26206 250392 26234
rect 249904 12374 249932 26206
rect 249984 24540 250036 24546
rect 249984 24482 250036 24488
rect 249892 12368 249944 12374
rect 249892 12310 249944 12316
rect 249800 11892 249852 11898
rect 249800 11834 249852 11840
rect 249996 480 250024 24482
rect 251192 3874 251220 35566
rect 251284 4554 251312 40035
rect 251836 26234 251864 40035
rect 252560 37868 252612 37874
rect 252560 37810 252612 37816
rect 251376 26206 251864 26234
rect 251376 6662 251404 26206
rect 251456 11892 251508 11898
rect 251456 11834 251508 11840
rect 251364 6656 251416 6662
rect 251364 6598 251416 6604
rect 251272 4548 251324 4554
rect 251272 4490 251324 4496
rect 251180 3868 251232 3874
rect 251180 3810 251232 3816
rect 251468 3482 251496 11834
rect 252572 6594 252600 37810
rect 252664 6866 252692 40035
rect 253584 37874 253612 40035
rect 253572 37868 253624 37874
rect 253572 37810 253624 37816
rect 254228 26234 254256 40035
rect 253952 26206 254256 26234
rect 252652 6860 252704 6866
rect 252652 6802 252704 6808
rect 252560 6588 252612 6594
rect 252560 6530 252612 6536
rect 253952 6526 253980 26206
rect 254216 12368 254268 12374
rect 254216 12310 254268 12316
rect 253940 6520 253992 6526
rect 253940 6462 253992 6468
rect 253480 6180 253532 6186
rect 253480 6122 253532 6128
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 251192 3454 251496 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3810
rect 253492 480 253520 6122
rect 248758 354 248870 480
rect 248616 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 12310
rect 255332 6390 255360 40174
rect 255792 40066 255820 40174
rect 263704 40174 264376 40202
rect 255424 6458 255452 40063
rect 255792 40038 256220 40066
rect 256712 40035 256980 40063
rect 257356 40035 257760 40063
rect 258092 40035 258560 40063
rect 258920 40035 259340 40063
rect 259748 40035 260120 40063
rect 260900 40035 261156 40063
rect 255504 19032 255556 19038
rect 255504 18974 255556 18980
rect 255516 16574 255544 18974
rect 255516 16546 255912 16574
rect 255412 6452 255464 6458
rect 255412 6394 255464 6400
rect 255320 6384 255372 6390
rect 255320 6326 255372 6332
rect 255884 480 255912 16546
rect 256712 6322 256740 40035
rect 257356 26234 257384 40035
rect 256804 26206 257384 26234
rect 256700 6316 256752 6322
rect 256700 6258 256752 6264
rect 256804 6254 256832 26206
rect 256884 21548 256936 21554
rect 256884 21490 256936 21496
rect 256792 6248 256844 6254
rect 256792 6190 256844 6196
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256896 354 256924 21490
rect 258092 5302 258120 40035
rect 258920 26234 258948 40035
rect 259748 35894 259776 40035
rect 261128 37874 261156 40035
rect 261220 40035 261680 40063
rect 262324 40035 262440 40063
rect 262876 40035 263220 40063
rect 261116 37868 261168 37874
rect 261116 37810 261168 37816
rect 259564 35866 259776 35894
rect 259460 34196 259512 34202
rect 259460 34138 259512 34144
rect 258184 26206 258948 26234
rect 258184 6186 258212 26206
rect 258172 6180 258224 6186
rect 258172 6122 258224 6128
rect 258080 5296 258132 5302
rect 258080 5238 258132 5244
rect 258264 4548 258316 4554
rect 258264 4490 258316 4496
rect 258276 480 258304 4490
rect 259472 480 259500 34138
rect 259564 7818 259592 35866
rect 261220 35358 261248 40035
rect 261208 35352 261260 35358
rect 261208 35294 261260 35300
rect 262220 28688 262272 28694
rect 262220 28630 262272 28636
rect 259644 28416 259696 28422
rect 259644 28358 259696 28364
rect 259656 16574 259684 28358
rect 262232 16574 262260 28630
rect 262324 21690 262352 40035
rect 262876 39930 262904 40035
rect 262784 39902 262904 39930
rect 262784 28762 262812 39902
rect 262864 37868 262916 37874
rect 262864 37810 262916 37816
rect 262772 28756 262824 28762
rect 262772 28698 262824 28704
rect 262312 21684 262364 21690
rect 262312 21626 262364 21632
rect 259656 16546 260696 16574
rect 262232 16546 262536 16574
rect 259552 7812 259604 7818
rect 259552 7754 259604 7760
rect 260668 480 260696 16546
rect 261760 6656 261812 6662
rect 261760 6598 261812 6604
rect 261772 480 261800 6598
rect 257038 354 257150 480
rect 256896 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 262876 15026 262904 37810
rect 263704 26234 263732 40174
rect 264348 40066 264376 40174
rect 267844 40174 268332 40202
rect 263612 26206 263732 26234
rect 263796 40035 264020 40063
rect 264348 40038 264800 40066
rect 265176 40035 265580 40063
rect 266360 40035 266492 40063
rect 262864 15020 262916 15026
rect 262864 14962 262916 14968
rect 263612 8158 263640 26206
rect 263796 23254 263824 40035
rect 265176 26234 265204 40035
rect 266360 37868 266412 37874
rect 266360 37810 266412 37816
rect 264992 26206 265204 26234
rect 263784 23248 263836 23254
rect 263784 23190 263836 23196
rect 263692 22908 263744 22914
rect 263692 22850 263744 22856
rect 263704 16574 263732 22850
rect 263704 16546 264192 16574
rect 263600 8152 263652 8158
rect 263600 8094 263652 8100
rect 264164 480 264192 16546
rect 264992 6730 265020 26206
rect 266372 12238 266400 37810
rect 266464 12306 266492 40035
rect 266832 40035 267140 40063
rect 266832 37874 266860 40035
rect 266820 37868 266872 37874
rect 266820 37810 266872 37816
rect 267844 35894 267872 40174
rect 268304 40066 268332 40174
rect 269132 40174 269896 40202
rect 267906 39794 267934 40049
rect 268304 40038 268700 40066
rect 267906 39766 267964 39794
rect 267752 35866 267872 35894
rect 266544 23180 266596 23186
rect 266544 23122 266596 23128
rect 266452 12300 266504 12306
rect 266452 12242 266504 12248
rect 266360 12232 266412 12238
rect 266360 12174 266412 12180
rect 265348 6860 265400 6866
rect 265348 6802 265400 6808
rect 264980 6724 265032 6730
rect 264980 6666 265032 6672
rect 265360 480 265388 6802
rect 266556 480 266584 23122
rect 267752 12170 267780 35866
rect 267832 27056 267884 27062
rect 267832 26998 267884 27004
rect 267740 12164 267792 12170
rect 267740 12106 267792 12112
rect 267844 6914 267872 26998
rect 267936 20398 267964 39766
rect 267924 20392 267976 20398
rect 267924 20334 267976 20340
rect 269132 12034 269160 40174
rect 269868 40066 269896 40174
rect 280172 40174 280844 40202
rect 269224 40035 269500 40063
rect 269868 40038 270280 40066
rect 270604 40035 271040 40063
rect 271432 40035 271820 40063
rect 272260 40035 272600 40063
rect 269224 12102 269252 40035
rect 270500 29776 270552 29782
rect 270500 29718 270552 29724
rect 269304 17672 269356 17678
rect 269304 17614 269356 17620
rect 269316 16574 269344 17614
rect 269316 16546 270080 16574
rect 269212 12096 269264 12102
rect 269212 12038 269264 12044
rect 269120 12028 269172 12034
rect 269120 11970 269172 11976
rect 267752 6886 267872 6914
rect 267752 480 267780 6886
rect 268844 6588 268896 6594
rect 268844 6530 268896 6536
rect 268856 480 268884 6530
rect 270052 480 270080 16546
rect 270512 6914 270540 29718
rect 270604 11966 270632 40035
rect 271432 26234 271460 40035
rect 272260 26234 272288 40035
rect 273260 31476 273312 31482
rect 273260 31418 273312 31424
rect 270696 26206 271460 26234
rect 271892 26206 272288 26234
rect 270592 11960 270644 11966
rect 270592 11902 270644 11908
rect 270696 11830 270724 26206
rect 271892 11898 271920 26206
rect 271880 11892 271932 11898
rect 271880 11834 271932 11840
rect 270684 11824 270736 11830
rect 270684 11766 270736 11772
rect 270512 6886 270816 6914
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 354 270816 6886
rect 272432 6520 272484 6526
rect 272432 6462 272484 6468
rect 272444 480 272472 6462
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 31418
rect 273364 11762 273392 40063
rect 273732 40035 274160 40063
rect 274940 40035 275232 40063
rect 275720 40035 275968 40063
rect 273732 27334 273760 40035
rect 275204 37330 275232 40035
rect 275192 37324 275244 37330
rect 275192 37266 275244 37272
rect 275940 32774 275968 40035
rect 276124 40035 276500 40063
rect 275928 32768 275980 32774
rect 275928 32710 275980 32716
rect 276124 30054 276152 40035
rect 277266 39794 277294 40049
rect 278060 40035 278360 40063
rect 278840 40035 279096 40063
rect 277228 39766 277294 39794
rect 277228 38214 277256 39766
rect 277216 38208 277268 38214
rect 277216 38150 277268 38156
rect 277400 36712 277452 36718
rect 277400 36654 277452 36660
rect 276112 30048 276164 30054
rect 276112 29990 276164 29996
rect 273720 27328 273772 27334
rect 273720 27270 273772 27276
rect 276020 24540 276072 24546
rect 276020 24482 276072 24488
rect 276032 16574 276060 24482
rect 277412 16574 277440 36654
rect 278332 34134 278360 40035
rect 279068 37670 279096 40035
rect 279252 40035 279640 40063
rect 279056 37664 279108 37670
rect 279056 37606 279108 37612
rect 278320 34128 278372 34134
rect 278320 34070 278372 34076
rect 279252 28626 279280 40035
rect 279240 28620 279292 28626
rect 279240 28562 279292 28568
rect 276032 16546 276704 16574
rect 277412 16546 278360 16574
rect 274824 13252 274876 13258
rect 274824 13194 274876 13200
rect 273352 11756 273404 11762
rect 273352 11698 273404 11704
rect 274836 480 274864 13194
rect 276020 6452 276072 6458
rect 276020 6394 276072 6400
rect 276032 480 276060 6394
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 280172 13734 280200 40174
rect 280816 40066 280844 40174
rect 287072 40174 287836 40202
rect 280264 40035 280420 40063
rect 280816 40038 281200 40066
rect 281552 40035 281980 40063
rect 282380 40035 282760 40063
rect 283116 40035 283540 40063
rect 284320 40035 284432 40063
rect 280264 18970 280292 40035
rect 280804 37664 280856 37670
rect 280804 37606 280856 37612
rect 280816 21826 280844 37606
rect 280804 21820 280856 21826
rect 280804 21762 280856 21768
rect 280252 18964 280304 18970
rect 280252 18906 280304 18912
rect 280712 14952 280764 14958
rect 280712 14894 280764 14900
rect 280160 13728 280212 13734
rect 280160 13670 280212 13676
rect 279516 6384 279568 6390
rect 279516 6326 279568 6332
rect 279528 480 279556 6326
rect 280724 480 280752 14894
rect 281552 13666 281580 40035
rect 282380 39930 282408 40035
rect 282104 39902 282408 39930
rect 282104 26234 282132 39902
rect 282184 38344 282236 38350
rect 282184 38286 282236 38292
rect 281644 26206 282132 26234
rect 281540 13660 281592 13666
rect 281540 13602 281592 13608
rect 281644 13598 281672 26206
rect 281724 14544 281776 14550
rect 281724 14486 281776 14492
rect 281632 13592 281684 13598
rect 281632 13534 281684 13540
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281736 354 281764 14486
rect 282196 13122 282224 38286
rect 283116 26234 283144 40035
rect 284300 37868 284352 37874
rect 284300 37810 284352 37816
rect 282932 26206 283144 26234
rect 282932 13530 282960 26206
rect 282920 13524 282972 13530
rect 282920 13466 282972 13472
rect 284312 13394 284340 37810
rect 284404 13462 284432 40035
rect 284772 40035 285100 40063
rect 285692 40035 285880 40063
rect 286244 40035 286640 40063
rect 284772 37874 284800 40035
rect 284760 37868 284812 37874
rect 284760 37810 284812 37816
rect 284484 20120 284536 20126
rect 284484 20062 284536 20068
rect 284496 16574 284524 20062
rect 284496 16546 284984 16574
rect 284392 13456 284444 13462
rect 284392 13398 284444 13404
rect 284300 13388 284352 13394
rect 284300 13330 284352 13336
rect 282184 13116 282236 13122
rect 282184 13058 282236 13064
rect 284300 8220 284352 8226
rect 284300 8162 284352 8168
rect 283104 6316 283156 6322
rect 283104 6258 283156 6264
rect 283116 480 283144 6258
rect 284312 480 284340 8162
rect 281878 354 281990 480
rect 281736 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 285692 13122 285720 40035
rect 286244 26234 286272 40035
rect 286324 38276 286376 38282
rect 286324 38218 286376 38224
rect 285784 26206 286272 26234
rect 285784 13326 285812 26206
rect 285772 13320 285824 13326
rect 285772 13262 285824 13268
rect 286336 13190 286364 38218
rect 287072 13190 287100 40174
rect 287808 40066 287836 40174
rect 298112 40174 298784 40202
rect 287164 40035 287420 40063
rect 287808 40038 288200 40066
rect 288636 40035 288980 40063
rect 289464 40035 289780 40063
rect 290108 40035 290560 40063
rect 291212 40035 291340 40063
rect 291764 40035 292120 40063
rect 292900 40035 293172 40063
rect 287164 13258 287192 40035
rect 288440 37868 288492 37874
rect 288440 37810 288492 37816
rect 288452 20126 288480 37810
rect 288636 26234 288664 40035
rect 289464 37874 289492 40035
rect 289452 37868 289504 37874
rect 289452 37810 289504 37816
rect 290108 35562 290136 40035
rect 290096 35556 290148 35562
rect 290096 35498 290148 35504
rect 288544 26206 288664 26234
rect 288544 23118 288572 26206
rect 288532 23112 288584 23118
rect 288532 23054 288584 23060
rect 288440 20120 288492 20126
rect 288440 20062 288492 20068
rect 288440 18760 288492 18766
rect 288440 18702 288492 18708
rect 288452 16574 288480 18702
rect 291212 17542 291240 40035
rect 291764 31346 291792 40035
rect 293144 37806 293172 40035
rect 293236 40035 293680 40063
rect 294156 40035 294460 40063
rect 294984 40035 295260 40063
rect 295628 40035 296040 40063
rect 296820 40035 297128 40063
rect 297600 40035 297864 40063
rect 293132 37800 293184 37806
rect 293132 37742 293184 37748
rect 291844 32836 291896 32842
rect 291844 32778 291896 32784
rect 291752 31340 291804 31346
rect 291752 31282 291804 31288
rect 291200 17536 291252 17542
rect 291200 17478 291252 17484
rect 288452 16546 289032 16574
rect 287152 13252 287204 13258
rect 287152 13194 287204 13200
rect 286324 13184 286376 13190
rect 286324 13126 286376 13132
rect 287060 13184 287112 13190
rect 287060 13126 287112 13132
rect 285680 13116 285732 13122
rect 285680 13058 285732 13064
rect 286600 6248 286652 6254
rect 286600 6190 286652 6196
rect 286612 480 286640 6190
rect 287796 3392 287848 3398
rect 287796 3334 287848 3340
rect 287808 480 287836 3334
rect 289004 480 289032 16546
rect 290188 5296 290240 5302
rect 290188 5238 290240 5244
rect 290200 480 290228 5238
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 291396 480 291424 3810
rect 291856 3398 291884 32778
rect 293236 26234 293264 40035
rect 294052 37868 294104 37874
rect 294052 37810 294104 37816
rect 293960 27396 294012 27402
rect 293960 27338 294012 27344
rect 292684 26206 293264 26234
rect 292580 25696 292632 25702
rect 292580 25638 292632 25644
rect 291844 3392 291896 3398
rect 291844 3334 291896 3340
rect 292592 480 292620 25638
rect 292684 16046 292712 26206
rect 293972 16574 294000 27338
rect 294064 25838 294092 37810
rect 294156 27266 294184 40035
rect 294984 37874 295012 40035
rect 294972 37868 295024 37874
rect 294972 37810 295024 37816
rect 295340 32632 295392 32638
rect 295340 32574 295392 32580
rect 294144 27260 294196 27266
rect 294144 27202 294196 27208
rect 294052 25832 294104 25838
rect 294052 25774 294104 25780
rect 294604 21888 294656 21894
rect 294604 21830 294656 21836
rect 293972 16546 294552 16574
rect 292672 16040 292724 16046
rect 292672 15982 292724 15988
rect 293684 6180 293736 6186
rect 293684 6122 293736 6128
rect 293696 480 293724 6122
rect 294524 3482 294552 16546
rect 294616 3874 294644 21830
rect 295352 6914 295380 32574
rect 295628 26234 295656 40035
rect 297100 38486 297128 40035
rect 297088 38480 297140 38486
rect 297088 38422 297140 38428
rect 295984 37800 296036 37806
rect 295984 37742 296036 37748
rect 295996 32638 296024 37742
rect 297836 36786 297864 40035
rect 297824 36780 297876 36786
rect 297824 36722 297876 36728
rect 295984 32632 296036 32638
rect 295984 32574 296036 32580
rect 295444 26206 295656 26234
rect 295444 14754 295472 26206
rect 295432 14748 295484 14754
rect 295432 14690 295484 14696
rect 298112 14618 298140 40174
rect 298756 40066 298784 40174
rect 299492 40174 300256 40202
rect 298204 40035 298380 40063
rect 298756 40038 299160 40066
rect 298204 14686 298232 40035
rect 298284 16448 298336 16454
rect 298284 16390 298336 16396
rect 298192 14680 298244 14686
rect 298192 14622 298244 14628
rect 298100 14612 298152 14618
rect 298100 14554 298152 14560
rect 297272 7812 297324 7818
rect 297272 7754 297324 7760
rect 295352 6886 295656 6914
rect 294604 3868 294656 3874
rect 294604 3810 294656 3816
rect 294524 3454 294920 3482
rect 294892 480 294920 3454
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 354 295656 6886
rect 297284 480 297312 7754
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298296 354 298324 16390
rect 299492 6662 299520 40174
rect 300228 40066 300256 40174
rect 303724 40174 304212 40202
rect 299584 40035 299920 40063
rect 300228 40038 300700 40066
rect 301056 40035 301480 40063
rect 299584 14550 299612 40035
rect 301056 26234 301084 40035
rect 300872 26206 301084 26234
rect 300768 15020 300820 15026
rect 300768 14962 300820 14968
rect 299572 14544 299624 14550
rect 299572 14486 299624 14492
rect 299664 7744 299716 7750
rect 299664 7686 299716 7692
rect 299480 6656 299532 6662
rect 299480 6598 299532 6604
rect 299676 480 299704 7686
rect 300780 480 300808 14962
rect 300872 6594 300900 26206
rect 300860 6588 300912 6594
rect 300860 6530 300912 6536
rect 302252 6526 302280 40063
rect 302620 40035 303040 40063
rect 302620 26234 302648 40035
rect 303620 35352 303672 35358
rect 303620 35294 303672 35300
rect 302344 26206 302648 26234
rect 302240 6520 302292 6526
rect 302240 6462 302292 6468
rect 302344 6458 302372 26206
rect 303160 7676 303212 7682
rect 303160 7618 303212 7624
rect 302332 6452 302384 6458
rect 302332 6394 302384 6400
rect 301964 2916 302016 2922
rect 301964 2858 302016 2864
rect 301976 480 302004 2858
rect 303172 480 303200 7618
rect 298438 354 298550 480
rect 298296 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303632 354 303660 35294
rect 303724 6322 303752 40174
rect 304184 40066 304212 40174
rect 327184 40174 327672 40202
rect 303816 6390 303844 40063
rect 304184 40038 304600 40066
rect 305012 40035 305400 40063
rect 305748 40035 306180 40063
rect 306576 40035 306960 40063
rect 307740 40035 308076 40063
rect 303804 6384 303856 6390
rect 303804 6326 303856 6332
rect 303712 6316 303764 6322
rect 303712 6258 303764 6264
rect 305012 6254 305040 40035
rect 305748 26234 305776 40035
rect 306576 26234 306604 40035
rect 307116 38208 307168 38214
rect 307116 38150 307168 38156
rect 307024 34264 307076 34270
rect 307024 34206 307076 34212
rect 305104 26206 305776 26234
rect 306392 26206 306604 26234
rect 305000 6248 305052 6254
rect 305000 6190 305052 6196
rect 305104 6186 305132 26206
rect 306392 21554 306420 26206
rect 306380 21548 306432 21554
rect 306380 21490 306432 21496
rect 306748 7608 306800 7614
rect 306748 7550 306800 7556
rect 305092 6180 305144 6186
rect 305092 6122 305144 6128
rect 305550 3360 305606 3369
rect 305550 3295 305606 3304
rect 305564 480 305592 3295
rect 306760 480 306788 7550
rect 307036 2922 307064 34206
rect 307128 20330 307156 38150
rect 308048 37874 308076 40035
rect 308140 40035 308520 40063
rect 309152 40035 309300 40063
rect 309612 40035 310080 40063
rect 310624 40035 310860 40063
rect 311640 40035 311848 40063
rect 308036 37868 308088 37874
rect 308036 37810 308088 37816
rect 308140 26234 308168 40035
rect 309152 27062 309180 40035
rect 309612 29782 309640 40035
rect 309784 37868 309836 37874
rect 309784 37810 309836 37816
rect 309600 29776 309652 29782
rect 309600 29718 309652 29724
rect 309796 28422 309824 37810
rect 310520 28756 310572 28762
rect 310520 28698 310572 28704
rect 309784 28416 309836 28422
rect 309784 28358 309836 28364
rect 309140 27056 309192 27062
rect 309140 26998 309192 27004
rect 307772 26206 308168 26234
rect 307772 22914 307800 26206
rect 309140 24268 309192 24274
rect 309140 24210 309192 24216
rect 307760 22908 307812 22914
rect 307760 22850 307812 22856
rect 307760 21684 307812 21690
rect 307760 21626 307812 21632
rect 307116 20324 307168 20330
rect 307116 20266 307168 20272
rect 307772 16574 307800 21626
rect 309152 16574 309180 24210
rect 310532 16574 310560 28698
rect 310624 18766 310652 40035
rect 311820 38418 311848 40035
rect 312004 40035 312420 40063
rect 311808 38412 311860 38418
rect 311808 38354 311860 38360
rect 312004 35358 312032 40035
rect 312544 38480 312596 38486
rect 312544 38422 312596 38428
rect 311992 35352 312044 35358
rect 311992 35294 312044 35300
rect 312556 21690 312584 38422
rect 313200 36718 313228 40063
rect 313568 40035 313980 40063
rect 314740 40035 315068 40063
rect 313188 36712 313240 36718
rect 313188 36654 313240 36660
rect 313280 33992 313332 33998
rect 313280 33934 313332 33940
rect 312544 21684 312596 21690
rect 312544 21626 312596 21632
rect 310612 18760 310664 18766
rect 310612 18702 310664 18708
rect 307772 16546 307984 16574
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 307024 2916 307076 2922
rect 307024 2858 307076 2864
rect 307956 480 307984 16546
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 309060 480 309088 3810
rect 304326 354 304438 480
rect 303632 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 313292 6914 313320 33934
rect 313568 26234 313596 40035
rect 315040 37330 315068 40035
rect 315132 40035 315520 40063
rect 316052 40035 316320 40063
rect 316696 40035 317100 40063
rect 317432 40035 317880 40063
rect 318260 40035 318660 40063
rect 318996 40035 319440 40063
rect 320220 40035 320312 40063
rect 315028 37324 315080 37330
rect 315028 37266 315080 37272
rect 315132 26234 315160 40035
rect 313384 26206 313596 26234
rect 314672 26206 315160 26234
rect 313384 8022 313412 26206
rect 314672 25702 314700 26206
rect 314660 25696 314712 25702
rect 314660 25638 314712 25644
rect 314660 23248 314712 23254
rect 314660 23190 314712 23196
rect 313372 8016 313424 8022
rect 313372 7958 313424 7964
rect 313292 6886 313872 6914
rect 312636 3936 312688 3942
rect 312636 3878 312688 3884
rect 312648 480 312676 3878
rect 313844 480 313872 6886
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 23190
rect 316052 7954 316080 40035
rect 316696 26234 316724 40035
rect 316144 26206 316724 26234
rect 316040 7948 316092 7954
rect 316040 7890 316092 7896
rect 316144 7886 316172 26206
rect 316224 21616 316276 21622
rect 316224 21558 316276 21564
rect 316236 16574 316264 21558
rect 316236 16546 317368 16574
rect 316132 7880 316184 7886
rect 316132 7822 316184 7828
rect 316224 4004 316276 4010
rect 316224 3946 316276 3952
rect 316236 480 316264 3946
rect 317340 480 317368 16546
rect 317432 7818 317460 40035
rect 318260 39386 318288 40035
rect 317984 39358 318288 39386
rect 317984 26234 318012 39358
rect 318064 37324 318116 37330
rect 318064 37266 318116 37272
rect 317524 26206 318012 26234
rect 317420 7812 317472 7818
rect 317420 7754 317472 7760
rect 317524 7750 317552 26206
rect 318076 15910 318104 37266
rect 318996 26234 319024 40035
rect 320180 37868 320232 37874
rect 320180 37810 320232 37816
rect 318812 26206 319024 26234
rect 318812 24274 318840 26206
rect 318800 24268 318852 24274
rect 318800 24210 318852 24216
rect 318064 15904 318116 15910
rect 318064 15846 318116 15852
rect 318524 8152 318576 8158
rect 318524 8094 318576 8100
rect 317512 7744 317564 7750
rect 317512 7686 317564 7692
rect 318536 480 318564 8094
rect 320192 7614 320220 37810
rect 320284 7682 320312 40035
rect 320744 40035 321020 40063
rect 321800 40035 322060 40063
rect 320744 37874 320772 40035
rect 322032 38214 322060 40035
rect 322124 40035 322580 40063
rect 323044 40035 323360 40063
rect 323780 40035 324120 40063
rect 324608 40035 324900 40063
rect 325680 40035 325832 40063
rect 322020 38208 322072 38214
rect 322020 38150 322072 38156
rect 320732 37868 320784 37874
rect 320732 37810 320784 37816
rect 320364 28552 320416 28558
rect 320364 28494 320416 28500
rect 320376 16574 320404 28494
rect 322124 26234 322152 40035
rect 323044 37874 323072 40035
rect 322204 37868 322256 37874
rect 322204 37810 322256 37816
rect 323032 37868 323084 37874
rect 323032 37810 323084 37816
rect 321572 26206 322152 26234
rect 320376 16546 320496 16574
rect 320272 7676 320324 7682
rect 320272 7618 320324 7624
rect 320180 7608 320232 7614
rect 320180 7550 320232 7556
rect 319720 4072 319772 4078
rect 319720 4014 319772 4020
rect 319732 480 319760 4014
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 321572 14482 321600 26206
rect 321560 14476 321612 14482
rect 321560 14418 321612 14424
rect 322216 8090 322244 37810
rect 323780 27130 323808 40035
rect 324608 38350 324636 40035
rect 324596 38344 324648 38350
rect 324596 38286 324648 38292
rect 324964 38344 325016 38350
rect 324964 38286 325016 38292
rect 323768 27124 323820 27130
rect 323768 27066 323820 27072
rect 324320 22976 324372 22982
rect 324320 22918 324372 22924
rect 322204 8084 322256 8090
rect 322204 8026 322256 8032
rect 322112 6724 322164 6730
rect 322112 6666 322164 6672
rect 322124 480 322152 6666
rect 323308 4140 323360 4146
rect 323308 4082 323360 4088
rect 323320 480 323348 4082
rect 324332 3210 324360 22918
rect 324412 12300 324464 12306
rect 324412 12242 324464 12248
rect 324424 3398 324452 12242
rect 324976 8226 325004 38286
rect 325700 37868 325752 37874
rect 325700 37810 325752 37816
rect 324964 8220 325016 8226
rect 324964 8162 325016 8168
rect 325712 3534 325740 37810
rect 325700 3528 325752 3534
rect 325700 3470 325752 3476
rect 325804 3466 325832 40035
rect 326172 40035 326480 40063
rect 326172 37874 326200 40035
rect 326160 37868 326212 37874
rect 326160 37810 326212 37816
rect 327080 36848 327132 36854
rect 327080 36790 327132 36796
rect 327092 3482 327120 36790
rect 327184 3670 327212 40174
rect 327644 40066 327672 40174
rect 333992 40174 334664 40202
rect 327246 39794 327274 40049
rect 327644 40038 328040 40066
rect 328472 40035 328800 40063
rect 329116 40035 329580 40063
rect 330036 40035 330360 40063
rect 330772 40035 331140 40063
rect 331508 40035 331940 40063
rect 332612 40035 332720 40063
rect 333072 40035 333500 40063
rect 327246 39766 327304 39794
rect 327172 3664 327224 3670
rect 327172 3606 327224 3612
rect 327276 3602 327304 39766
rect 328472 3738 328500 40035
rect 328736 38072 328788 38078
rect 328736 38014 328788 38020
rect 328748 37874 328776 38014
rect 328736 37868 328788 37874
rect 328736 37810 328788 37816
rect 329116 26234 329144 40035
rect 330036 38282 330064 40035
rect 330772 39352 330800 40035
rect 330404 39324 330800 39352
rect 330024 38276 330076 38282
rect 330024 38218 330076 38224
rect 330404 35494 330432 39324
rect 330576 38276 330628 38282
rect 330576 38218 330628 38224
rect 330484 38072 330536 38078
rect 330484 38014 330536 38020
rect 330392 35488 330444 35494
rect 330392 35430 330444 35436
rect 328564 26206 329144 26234
rect 328564 3806 328592 26206
rect 330496 18902 330524 38014
rect 330588 25974 330616 38218
rect 331220 27192 331272 27198
rect 331220 27134 331272 27140
rect 330576 25968 330628 25974
rect 330576 25910 330628 25916
rect 330484 18896 330536 18902
rect 330484 18838 330536 18844
rect 328736 12232 328788 12238
rect 328736 12174 328788 12180
rect 328552 3800 328604 3806
rect 328552 3742 328604 3748
rect 328460 3732 328512 3738
rect 328460 3674 328512 3680
rect 327264 3596 327316 3602
rect 327264 3538 327316 3544
rect 325792 3460 325844 3466
rect 325792 3402 325844 3408
rect 326804 3460 326856 3466
rect 327092 3454 328040 3482
rect 326804 3402 326856 3408
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 326816 480 326844 3402
rect 328012 480 328040 3454
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 12174
rect 330392 3528 330444 3534
rect 330392 3470 330444 3476
rect 330404 480 330432 3470
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 27134
rect 331508 26234 331536 40035
rect 332612 38078 332640 40035
rect 332600 38072 332652 38078
rect 332600 38014 332652 38020
rect 331864 37868 331916 37874
rect 331864 37810 331916 37816
rect 331324 26206 331536 26234
rect 331324 14822 331352 26206
rect 331876 16250 331904 37810
rect 333072 28490 333100 40035
rect 333060 28484 333112 28490
rect 333060 28426 333112 28432
rect 333992 24410 334020 40174
rect 334636 40066 334664 40174
rect 345032 40174 345612 40202
rect 334084 40035 334280 40063
rect 334636 40038 335060 40066
rect 335464 40035 335840 40063
rect 336292 40035 336620 40063
rect 337028 40035 337400 40063
rect 333980 24404 334032 24410
rect 333980 24346 334032 24352
rect 332600 20392 332652 20398
rect 332600 20334 332652 20340
rect 332612 16574 332640 20334
rect 332612 16546 332732 16574
rect 331864 16244 331916 16250
rect 331864 16186 331916 16192
rect 331312 14816 331364 14822
rect 331312 14758 331364 14764
rect 332704 480 332732 16546
rect 334084 15978 334112 40035
rect 335360 38072 335412 38078
rect 335360 38014 335412 38020
rect 334164 29844 334216 29850
rect 334164 29786 334216 29792
rect 334176 16574 334204 29786
rect 334176 16546 334664 16574
rect 334072 15972 334124 15978
rect 334072 15914 334124 15920
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 333900 480 333928 3538
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335372 16182 335400 38014
rect 335360 16176 335412 16182
rect 335360 16118 335412 16124
rect 335464 16114 335492 40035
rect 336292 38078 336320 40035
rect 336280 38072 336332 38078
rect 336280 38014 336332 38020
rect 337028 26234 337056 40035
rect 338166 39794 338194 40049
rect 336752 26206 337056 26234
rect 338132 39766 338194 39794
rect 338500 40035 338960 40063
rect 339512 40035 339740 40063
rect 340064 40035 340520 40063
rect 340892 40035 341300 40063
rect 341628 40035 342100 40063
rect 342456 40035 342860 40063
rect 343640 40035 343680 40063
rect 336752 23050 336780 26206
rect 336740 23044 336792 23050
rect 336740 22986 336792 22992
rect 338132 16318 338160 39766
rect 338500 26234 338528 40035
rect 339512 29918 339540 40035
rect 340064 34066 340092 40035
rect 340892 38078 340920 40035
rect 341628 39930 341656 40035
rect 340984 39902 341656 39930
rect 340144 38072 340196 38078
rect 340144 38014 340196 38020
rect 340880 38072 340932 38078
rect 340880 38014 340932 38020
rect 340052 34060 340104 34066
rect 340052 34002 340104 34008
rect 339500 29912 339552 29918
rect 339500 29854 339552 29860
rect 338224 26206 338528 26234
rect 338224 25906 338252 26206
rect 338212 25900 338264 25906
rect 338212 25842 338264 25848
rect 338212 20188 338264 20194
rect 338212 20130 338264 20136
rect 338224 16574 338252 20130
rect 340156 17610 340184 38014
rect 340984 31414 341012 39902
rect 341064 38072 341116 38078
rect 341064 38014 341116 38020
rect 340972 31408 341024 31414
rect 340972 31350 341024 31356
rect 341076 26234 341104 38014
rect 342456 26234 342484 40035
rect 343652 38570 343680 40035
rect 343560 38542 343680 38570
rect 344020 40035 344420 40063
rect 342904 38140 342956 38146
rect 342904 38082 342956 38088
rect 340892 26206 341104 26234
rect 342272 26206 342484 26234
rect 340144 17604 340196 17610
rect 340144 17546 340196 17552
rect 338224 16546 338712 16574
rect 338120 16312 338172 16318
rect 338120 16254 338172 16260
rect 335452 16108 335504 16114
rect 335452 16050 335504 16056
rect 336280 12164 336332 12170
rect 336280 12106 336332 12112
rect 336292 480 336320 12106
rect 337476 3664 337528 3670
rect 337476 3606 337528 3612
rect 337488 480 337516 3606
rect 338684 480 338712 16546
rect 339500 12096 339552 12102
rect 339500 12038 339552 12044
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 12038
rect 340892 3210 340920 26206
rect 342272 21758 342300 26206
rect 342260 21752 342312 21758
rect 342260 21694 342312 21700
rect 340972 17468 341024 17474
rect 340972 17410 341024 17416
rect 340984 3398 341012 17410
rect 342916 15978 342944 38082
rect 343560 36922 343588 38542
rect 343548 36916 343600 36922
rect 343548 36858 343600 36864
rect 344020 26234 344048 40035
rect 345032 32706 345060 40174
rect 345584 40066 345612 40174
rect 351932 40174 352696 40202
rect 345124 40035 345200 40063
rect 345584 40038 345980 40066
rect 346412 40035 346760 40063
rect 347148 40035 347560 40063
rect 347884 40035 348320 40063
rect 348804 40035 349100 40063
rect 349540 40035 349880 40063
rect 350552 40035 350660 40063
rect 351012 40035 351440 40063
rect 345020 32700 345072 32706
rect 345020 32642 345072 32648
rect 345020 31272 345072 31278
rect 345020 31214 345072 31220
rect 343744 26206 344048 26234
rect 343744 16386 343772 26206
rect 343732 16380 343784 16386
rect 343732 16322 343784 16328
rect 342904 15972 342956 15978
rect 342904 15914 342956 15920
rect 342904 12028 342956 12034
rect 342904 11970 342956 11976
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 11970
rect 345032 6914 345060 31214
rect 345124 14890 345152 40035
rect 346412 20262 346440 40035
rect 347148 26234 347176 40035
rect 347884 29986 347912 40035
rect 348804 38282 348832 40035
rect 348792 38276 348844 38282
rect 348792 38218 348844 38224
rect 348424 37868 348476 37874
rect 348424 37810 348476 37816
rect 347872 29980 347924 29986
rect 347872 29922 347924 29928
rect 346504 26206 347176 26234
rect 346504 24478 346532 26206
rect 346492 24472 346544 24478
rect 346492 24414 346544 24420
rect 346400 20256 346452 20262
rect 346400 20198 346452 20204
rect 348436 19038 348464 37810
rect 349540 35630 349568 40035
rect 349804 38412 349856 38418
rect 349804 38354 349856 38360
rect 349528 35624 349580 35630
rect 349528 35566 349580 35572
rect 349160 35420 349212 35426
rect 349160 35362 349212 35368
rect 348424 19032 348476 19038
rect 348424 18974 348476 18980
rect 345112 14884 345164 14890
rect 345112 14826 345164 14832
rect 346952 11960 347004 11966
rect 346952 11902 347004 11908
rect 345032 6886 345336 6914
rect 344560 3732 344612 3738
rect 344560 3674 344612 3680
rect 344572 480 344600 3674
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 6886
rect 346964 480 346992 11902
rect 348056 3800 348108 3806
rect 348056 3742 348108 3748
rect 348068 480 348096 3742
rect 349172 3210 349200 35362
rect 349816 11830 349844 38354
rect 350552 37874 350580 40035
rect 350540 37868 350592 37874
rect 350540 37810 350592 37816
rect 351012 34202 351040 40035
rect 351000 34196 351052 34202
rect 351000 34138 351052 34144
rect 351932 23186 351960 40174
rect 352668 40066 352696 40174
rect 357452 40174 358124 40202
rect 352024 40035 352240 40063
rect 352668 40038 353020 40066
rect 353312 40035 353800 40063
rect 354140 40035 354580 40063
rect 355060 40035 355360 40063
rect 352024 28694 352052 40035
rect 352012 28688 352064 28694
rect 352012 28630 352064 28636
rect 351920 23180 351972 23186
rect 351920 23122 351972 23128
rect 351920 18828 351972 18834
rect 351920 18770 351972 18776
rect 351932 16574 351960 18770
rect 353312 17678 353340 40035
rect 354140 38842 354168 40035
rect 353864 38814 354168 38842
rect 353864 31482 353892 38814
rect 355060 37330 355088 40035
rect 356126 39794 356154 40049
rect 356624 40035 356920 40063
rect 356126 39766 356192 39794
rect 353944 37324 353996 37330
rect 353944 37266 353996 37272
rect 355048 37324 355100 37330
rect 355048 37266 355100 37272
rect 353852 31476 353904 31482
rect 353852 31418 353904 31424
rect 353956 24546 353984 37266
rect 353944 24540 353996 24546
rect 353944 24482 353996 24488
rect 353300 17672 353352 17678
rect 353300 17614 353352 17620
rect 351932 16546 352880 16574
rect 349252 11824 349304 11830
rect 349252 11766 349304 11772
rect 349804 11824 349856 11830
rect 349804 11766 349856 11772
rect 349264 3398 349292 11766
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 351644 3392 351696 3398
rect 351644 3334 351696 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 351656 480 351684 3334
rect 352852 480 352880 16546
rect 356164 14958 356192 39766
rect 356624 38350 356652 40035
rect 356612 38344 356664 38350
rect 356612 38286 356664 38292
rect 356704 38004 356756 38010
rect 356704 37946 356756 37952
rect 356716 27402 356744 37946
rect 356704 27396 356756 27402
rect 356704 27338 356756 27344
rect 357452 21894 357480 40174
rect 358096 40066 358124 40174
rect 362972 40174 363552 40202
rect 357544 40035 357700 40063
rect 358096 40038 358480 40066
rect 358924 40035 359260 40063
rect 359660 40035 360040 40063
rect 360396 40035 360800 40063
rect 361580 40035 361620 40063
rect 357544 32842 357572 40035
rect 358924 38010 358952 40035
rect 358912 38004 358964 38010
rect 358912 37946 358964 37952
rect 357532 32836 357584 32842
rect 357532 32778 357584 32784
rect 359660 26234 359688 40035
rect 360396 34270 360424 40035
rect 360844 37868 360896 37874
rect 360844 37810 360896 37816
rect 360384 34264 360436 34270
rect 360384 34206 360436 34212
rect 360200 27328 360252 27334
rect 360200 27270 360252 27276
rect 358924 26206 359688 26234
rect 357440 21888 357492 21894
rect 357440 21830 357492 21836
rect 358924 16454 358952 26206
rect 358912 16448 358964 16454
rect 358912 16390 358964 16396
rect 356152 14952 356204 14958
rect 356152 14894 356204 14900
rect 353576 11892 353628 11898
rect 353576 11834 353628 11840
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 11834
rect 357532 11756 357584 11762
rect 357532 11698 357584 11704
rect 356336 9580 356388 9586
rect 356336 9522 356388 9528
rect 355232 3324 355284 3330
rect 355232 3266 355284 3272
rect 355244 480 355272 3266
rect 356348 480 356376 9522
rect 357544 480 357572 11698
rect 359924 9512 359976 9518
rect 359924 9454 359976 9460
rect 358728 3120 358780 3126
rect 358728 3062 358780 3068
rect 358740 480 358768 3062
rect 359936 480 359964 9454
rect 360212 6914 360240 27270
rect 360856 11762 360884 37810
rect 360844 11756 360896 11762
rect 360844 11698 360896 11704
rect 360212 6886 361160 6914
rect 361132 480 361160 6886
rect 361592 3369 361620 40035
rect 361960 40035 362360 40063
rect 361960 26234 361988 40035
rect 361684 26206 361988 26234
rect 361684 3874 361712 26206
rect 362972 4010 363000 40174
rect 363524 40066 363552 40174
rect 404372 40174 404952 40202
rect 363064 40035 363160 40063
rect 363524 40038 363940 40066
rect 364444 40035 364720 40063
rect 365088 40035 365500 40063
rect 365916 40035 366280 40063
rect 366744 40035 367060 40063
rect 367388 40035 367860 40063
rect 362960 4004 363012 4010
rect 362960 3946 363012 3952
rect 363064 3942 363092 40035
rect 364340 36984 364392 36990
rect 364340 36926 364392 36932
rect 363512 9444 363564 9450
rect 363512 9386 363564 9392
rect 363052 3936 363104 3942
rect 363052 3878 363104 3884
rect 361672 3868 361724 3874
rect 361672 3810 361724 3816
rect 362316 3868 362368 3874
rect 362316 3810 362368 3816
rect 361578 3360 361634 3369
rect 361578 3295 361634 3304
rect 362328 480 362356 3810
rect 363524 480 363552 9386
rect 364352 3482 364380 36926
rect 364444 4078 364472 40035
rect 365088 26234 365116 40035
rect 365720 38004 365772 38010
rect 365720 37946 365772 37952
rect 364536 26206 365116 26234
rect 364536 4146 364564 26206
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 364432 4072 364484 4078
rect 364432 4014 364484 4020
rect 365732 3534 365760 37946
rect 365916 26234 365944 40035
rect 366744 38010 366772 40035
rect 366732 38004 366784 38010
rect 366732 37946 366784 37952
rect 367388 35894 367416 40035
rect 368626 39794 368654 40049
rect 365824 26206 365944 26234
rect 367112 35866 367416 35894
rect 368584 39766 368654 39794
rect 369136 40035 369420 40063
rect 369872 40035 370200 40063
rect 370516 40035 370980 40063
rect 371252 40035 371740 40063
rect 372172 40035 372520 40063
rect 372908 40035 373300 40063
rect 365824 16574 365852 26206
rect 365824 16546 365944 16574
rect 365720 3528 365772 3534
rect 364352 3454 364656 3482
rect 365720 3470 365772 3476
rect 364628 480 364656 3454
rect 365812 3460 365864 3466
rect 365812 3402 365864 3408
rect 365824 480 365852 3402
rect 365916 3398 365944 16546
rect 367008 9376 367060 9382
rect 367008 9318 367060 9324
rect 365904 3392 365956 3398
rect 365904 3334 365956 3340
rect 367020 480 367048 9318
rect 367112 3602 367140 35866
rect 367192 32768 367244 32774
rect 367192 32710 367244 32716
rect 367204 16574 367232 32710
rect 367204 16546 367784 16574
rect 367100 3596 367152 3602
rect 367100 3538 367152 3544
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 368584 3670 368612 39766
rect 369136 38078 369164 40035
rect 369124 38072 369176 38078
rect 369124 38014 369176 38020
rect 369872 3738 369900 40035
rect 370516 26234 370544 40035
rect 369964 26206 370544 26234
rect 369964 3806 369992 26206
rect 370596 9308 370648 9314
rect 370596 9250 370648 9256
rect 369952 3800 370004 3806
rect 369952 3742 370004 3748
rect 369860 3732 369912 3738
rect 369860 3674 369912 3680
rect 368572 3664 368624 3670
rect 368572 3606 368624 3612
rect 369400 3188 369452 3194
rect 369400 3130 369452 3136
rect 369412 480 369440 3130
rect 370608 480 370636 9250
rect 371252 3330 371280 40035
rect 372172 35894 372200 40035
rect 371344 35866 372200 35894
rect 371240 3324 371292 3330
rect 371240 3266 371292 3272
rect 371344 3262 371372 35866
rect 371424 30048 371476 30054
rect 371424 29990 371476 29996
rect 371332 3256 371384 3262
rect 371332 3198 371384 3204
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371436 354 371464 29990
rect 372908 26234 372936 40035
rect 374066 39794 374094 40049
rect 372632 26206 372936 26234
rect 374012 39766 374094 39794
rect 374472 40035 374860 40063
rect 375484 40035 375640 40063
rect 376036 40035 376420 40063
rect 376864 40035 377200 40063
rect 377508 40035 377980 40063
rect 378428 40035 378780 40063
rect 372632 3126 372660 26206
rect 374012 3874 374040 39766
rect 374472 26234 374500 40035
rect 375380 38276 375432 38282
rect 375380 38218 375432 38224
rect 374104 26206 374500 26234
rect 374104 11778 374132 26206
rect 374184 20324 374236 20330
rect 374184 20266 374236 20272
rect 374196 16574 374224 20266
rect 374196 16546 375328 16574
rect 374104 11750 374224 11778
rect 374092 9240 374144 9246
rect 374092 9182 374144 9188
rect 374000 3868 374052 3874
rect 374000 3810 374052 3816
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372620 3120 372672 3126
rect 372620 3062 372672 3068
rect 372908 480 372936 3674
rect 374104 480 374132 9182
rect 374196 3466 374224 11750
rect 374184 3460 374236 3466
rect 374184 3402 374236 3408
rect 375300 480 375328 16546
rect 375392 1306 375420 38218
rect 375484 3194 375512 40035
rect 376036 26234 376064 40035
rect 376864 38282 376892 40035
rect 376852 38276 376904 38282
rect 376852 38218 376904 38224
rect 377508 26234 377536 40035
rect 378428 35894 378456 40035
rect 375576 26206 376064 26234
rect 376956 26206 377536 26234
rect 378152 35866 378456 35894
rect 375576 3738 375604 26206
rect 375564 3732 375616 3738
rect 375564 3674 375616 3680
rect 376956 3330 376984 26206
rect 377680 9172 377732 9178
rect 377680 9114 377732 9120
rect 376944 3324 376996 3330
rect 376944 3266 376996 3272
rect 375472 3188 375524 3194
rect 375472 3130 375524 3136
rect 375392 1278 376064 1306
rect 371670 354 371782 480
rect 371436 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 1278
rect 377692 480 377720 9114
rect 378152 2990 378180 35866
rect 378232 34128 378284 34134
rect 378232 34070 378284 34076
rect 378244 16574 378272 34070
rect 378244 16546 378456 16574
rect 378140 2984 378192 2990
rect 378140 2926 378192 2932
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379532 3874 379560 40063
rect 379900 40035 380340 40063
rect 380912 40035 381120 40063
rect 381556 40035 381900 40063
rect 382680 40035 382872 40063
rect 379900 26234 379928 40035
rect 379624 26206 379928 26234
rect 379520 3868 379572 3874
rect 379520 3810 379572 3816
rect 379624 3806 379652 26206
rect 379612 3800 379664 3806
rect 379612 3742 379664 3748
rect 380912 3738 380940 40035
rect 381556 26234 381584 40035
rect 382844 38078 382872 40035
rect 383028 40035 383480 40063
rect 383856 40035 384260 40063
rect 385020 40035 385172 40063
rect 382832 38072 382884 38078
rect 382832 38014 382884 38020
rect 383028 26234 383056 40035
rect 383856 26234 383884 40035
rect 385040 38004 385092 38010
rect 385040 37946 385092 37952
rect 381004 26206 381584 26234
rect 382292 26206 383056 26234
rect 383672 26206 383884 26234
rect 381004 9246 381032 26206
rect 382292 9314 382320 26206
rect 382372 21820 382424 21826
rect 382372 21762 382424 21768
rect 382280 9308 382332 9314
rect 382280 9250 382332 9256
rect 380992 9240 381044 9246
rect 380992 9182 381044 9188
rect 381176 9104 381228 9110
rect 381176 9046 381228 9052
rect 380900 3732 380952 3738
rect 380900 3674 380952 3680
rect 379980 3324 380032 3330
rect 379980 3266 380032 3272
rect 379992 480 380020 3266
rect 381188 480 381216 9046
rect 382384 480 382412 21762
rect 383672 11966 383700 26206
rect 383660 11960 383712 11966
rect 383660 11902 383712 11908
rect 384764 9036 384816 9042
rect 384764 8978 384816 8984
rect 383568 2984 383620 2990
rect 383568 2926 383620 2932
rect 383580 480 383608 2926
rect 384776 480 384804 8978
rect 385052 3942 385080 37946
rect 385040 3936 385092 3942
rect 385040 3878 385092 3884
rect 385144 3670 385172 40035
rect 385512 40035 385800 40063
rect 386432 40035 386560 40063
rect 386892 40035 387340 40063
rect 387812 40035 388120 40063
rect 388548 40035 388920 40063
rect 389284 40035 389700 40063
rect 390112 40035 390480 40063
rect 390848 40035 391260 40063
rect 391952 40035 392040 40063
rect 392820 40035 393084 40063
rect 385512 38010 385540 40035
rect 385500 38004 385552 38010
rect 385500 37946 385552 37952
rect 385224 28620 385276 28626
rect 385224 28562 385276 28568
rect 385236 16574 385264 28562
rect 385236 16546 386000 16574
rect 385132 3664 385184 3670
rect 385132 3606 385184 3612
rect 385972 480 386000 16546
rect 386432 3602 386460 40035
rect 386892 26234 386920 40035
rect 386524 26206 386920 26234
rect 386420 3596 386472 3602
rect 386420 3538 386472 3544
rect 386524 3466 386552 26206
rect 387156 3868 387208 3874
rect 387156 3810 387208 3816
rect 386512 3460 386564 3466
rect 386512 3402 386564 3408
rect 387168 480 387196 3810
rect 387812 3262 387840 40035
rect 388548 26234 388576 40035
rect 389180 38004 389232 38010
rect 389180 37946 389232 37952
rect 387904 26206 388576 26234
rect 387904 3330 387932 26206
rect 388260 8968 388312 8974
rect 388260 8910 388312 8916
rect 387892 3324 387944 3330
rect 387892 3266 387944 3272
rect 387800 3256 387852 3262
rect 387800 3198 387852 3204
rect 388272 480 388300 8910
rect 389192 4146 389220 37946
rect 389180 4140 389232 4146
rect 389180 4082 389232 4088
rect 389284 3398 389312 40035
rect 390112 38010 390140 40035
rect 390100 38004 390152 38010
rect 390100 37946 390152 37952
rect 390848 26234 390876 40035
rect 390572 26206 390876 26234
rect 389364 18964 389416 18970
rect 389364 18906 389416 18912
rect 389376 16574 389404 18906
rect 389376 16546 389496 16574
rect 389272 3392 389324 3398
rect 389272 3334 389324 3340
rect 389468 480 389496 16546
rect 390572 4078 390600 26206
rect 390652 25764 390704 25770
rect 390652 25706 390704 25712
rect 390560 4072 390612 4078
rect 390560 4014 390612 4020
rect 390560 3800 390612 3806
rect 390560 3742 390612 3748
rect 390572 1986 390600 3742
rect 390664 3534 390692 25706
rect 391952 4010 391980 40035
rect 393056 38282 393084 40035
rect 393332 40035 393600 40063
rect 394400 40035 394648 40063
rect 393044 38276 393096 38282
rect 393044 38218 393096 38224
rect 392584 38072 392636 38078
rect 392584 38014 392636 38020
rect 392492 13728 392544 13734
rect 392492 13670 392544 13676
rect 392504 6914 392532 13670
rect 392596 8974 392624 38014
rect 392584 8968 392636 8974
rect 392584 8910 392636 8916
rect 392504 6886 392624 6914
rect 391940 4004 391992 4010
rect 391940 3946 391992 3952
rect 392032 3936 392084 3942
rect 392032 3878 392084 3884
rect 392044 3602 392072 3878
rect 392032 3596 392084 3602
rect 392032 3538 392084 3544
rect 390652 3528 390704 3534
rect 390652 3470 390704 3476
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390572 1958 390692 1986
rect 390664 480 390692 1958
rect 391860 480 391888 3470
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 6886
rect 393332 3942 393360 40035
rect 394620 38146 394648 40035
rect 394804 40035 395180 40063
rect 394608 38140 394660 38146
rect 394608 38082 394660 38088
rect 393964 37936 394016 37942
rect 393964 37878 394016 37884
rect 393976 12034 394004 37878
rect 394804 35894 394832 40035
rect 395946 39794 395974 40049
rect 395908 39766 395974 39794
rect 396276 40035 396740 40063
rect 397520 40035 397776 40063
rect 395908 38078 395936 39766
rect 395896 38072 395948 38078
rect 395896 38014 395948 38020
rect 394712 35866 394832 35894
rect 393964 12028 394016 12034
rect 393964 11970 394016 11976
rect 393320 3936 393372 3942
rect 393320 3878 393372 3884
rect 394712 3874 394740 35866
rect 394792 32564 394844 32570
rect 394792 32506 394844 32512
rect 394804 16574 394832 32506
rect 396276 26234 396304 40035
rect 397748 38010 397776 40035
rect 397932 40035 398280 40063
rect 399080 40035 399340 40063
rect 397736 38004 397788 38010
rect 397736 37946 397788 37952
rect 397932 26234 397960 40035
rect 399312 37942 399340 40035
rect 399404 40035 399860 40063
rect 400232 40035 400620 40063
rect 401060 40035 401400 40063
rect 401796 40035 402180 40063
rect 402960 40035 403204 40063
rect 399300 37936 399352 37942
rect 399300 37878 399352 37884
rect 399404 26234 399432 40035
rect 396092 26206 396304 26234
rect 397472 26206 397960 26234
rect 398852 26206 399432 26234
rect 394804 16546 395384 16574
rect 394700 3868 394752 3874
rect 394700 3810 394752 3816
rect 394240 3732 394292 3738
rect 394240 3674 394292 3680
rect 394252 480 394280 3674
rect 395356 480 395384 16546
rect 396092 3806 396120 26206
rect 396172 13660 396224 13666
rect 396172 13602 396224 13608
rect 396080 3800 396132 3806
rect 396080 3742 396132 3748
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396184 354 396212 13602
rect 397472 3738 397500 26206
rect 397736 9240 397788 9246
rect 397736 9182 397788 9188
rect 397460 3732 397512 3738
rect 397460 3674 397512 3680
rect 397748 480 397776 9182
rect 398852 3369 398880 26206
rect 398932 24336 398984 24342
rect 398932 24278 398984 24284
rect 398838 3360 398894 3369
rect 398838 3295 398894 3304
rect 398944 480 398972 24278
rect 400128 13592 400180 13598
rect 400128 13534 400180 13540
rect 400140 480 400168 13534
rect 400232 9246 400260 40035
rect 401060 26234 401088 40035
rect 401796 26234 401824 40035
rect 402980 35896 403032 35902
rect 402980 35838 403032 35844
rect 400324 26206 401088 26234
rect 401612 26206 401824 26234
rect 400220 9240 400272 9246
rect 400220 9182 400272 9188
rect 400324 9178 400352 26206
rect 400312 9172 400364 9178
rect 400312 9114 400364 9120
rect 401612 9110 401640 26206
rect 401692 21480 401744 21486
rect 401692 21422 401744 21428
rect 401704 16574 401732 21422
rect 401704 16546 402560 16574
rect 401600 9104 401652 9110
rect 401600 9046 401652 9052
rect 401324 8968 401376 8974
rect 401324 8910 401376 8916
rect 401336 480 401364 8910
rect 402532 480 402560 16546
rect 402992 8974 403020 35838
rect 403176 26234 403204 40035
rect 403360 40035 403740 40063
rect 403360 35902 403388 40035
rect 403348 35896 403400 35902
rect 403348 35838 403400 35844
rect 403084 26206 403204 26234
rect 403084 9042 403112 26206
rect 404372 13530 404400 40174
rect 404924 40066 404952 40174
rect 412744 40174 413508 40202
rect 404464 40035 404540 40063
rect 404924 40038 405320 40066
rect 405752 40035 406100 40063
rect 406488 40035 406880 40063
rect 407316 40035 407660 40063
rect 408144 40035 408440 40063
rect 408788 40035 409220 40063
rect 409892 40035 410000 40063
rect 410352 40035 410780 40063
rect 411560 40035 411852 40063
rect 404464 28490 404492 40035
rect 405752 29918 405780 40035
rect 405740 29912 405792 29918
rect 405740 29854 405792 29860
rect 404452 28484 404504 28490
rect 404452 28426 404504 28432
rect 405740 28348 405792 28354
rect 405740 28290 405792 28296
rect 403624 13524 403676 13530
rect 403624 13466 403676 13472
rect 404360 13524 404412 13530
rect 404360 13466 404412 13472
rect 403072 9036 403124 9042
rect 403072 8978 403124 8984
rect 402980 8968 403032 8974
rect 402980 8910 403032 8916
rect 403636 480 403664 13466
rect 404820 9308 404872 9314
rect 404820 9250 404872 9256
rect 404832 480 404860 9250
rect 405752 6914 405780 28290
rect 406488 26234 406516 40035
rect 407120 35896 407172 35902
rect 407120 35838 407172 35844
rect 405844 26206 406516 26234
rect 405844 11898 405872 26206
rect 407132 18834 407160 35838
rect 407316 26234 407344 40035
rect 408144 35902 408172 40035
rect 408132 35896 408184 35902
rect 408132 35838 408184 35844
rect 408788 33998 408816 40035
rect 408776 33992 408828 33998
rect 408776 33934 408828 33940
rect 407224 26206 407344 26234
rect 407224 22982 407252 26206
rect 407212 22976 407264 22982
rect 407212 22918 407264 22924
rect 408500 22840 408552 22846
rect 408500 22782 408552 22788
rect 407120 18828 407172 18834
rect 407120 18770 407172 18776
rect 408512 16574 408540 22782
rect 409892 20194 409920 40035
rect 410352 26234 410380 40035
rect 411824 38350 411852 40035
rect 411916 40035 412340 40063
rect 411812 38344 411864 38350
rect 411812 38286 411864 38292
rect 411916 26234 411944 40035
rect 412640 36576 412692 36582
rect 412640 36518 412692 36524
rect 409984 26206 410380 26234
rect 411272 26206 411944 26234
rect 409984 21486 410012 26206
rect 409972 21480 410024 21486
rect 409972 21422 410024 21428
rect 409880 20188 409932 20194
rect 409880 20130 409932 20136
rect 408512 16546 409184 16574
rect 407120 13456 407172 13462
rect 407120 13398 407172 13404
rect 405832 11892 405884 11898
rect 405832 11834 405884 11840
rect 405752 6886 406056 6914
rect 406028 480 406056 6886
rect 407028 3664 407080 3670
rect 407028 3606 407080 3612
rect 407040 3194 407068 3606
rect 407132 3482 407160 13398
rect 407212 11960 407264 11966
rect 407212 11902 407264 11908
rect 407224 3670 407252 11902
rect 407212 3664 407264 3670
rect 407212 3606 407264 3612
rect 408408 3664 408460 3670
rect 408408 3606 408460 3612
rect 407132 3454 407252 3482
rect 407028 3188 407080 3194
rect 407028 3130 407080 3136
rect 407224 480 407252 3454
rect 408420 480 408448 3606
rect 396510 354 396622 480
rect 396184 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 411272 13394 411300 26206
rect 410800 13388 410852 13394
rect 410800 13330 410852 13336
rect 411260 13388 411312 13394
rect 411260 13330 411312 13336
rect 410812 480 410840 13330
rect 411904 3188 411956 3194
rect 411904 3130 411956 3136
rect 411916 480 411944 3130
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 36518
rect 412744 24342 412772 40174
rect 413480 40066 413508 40174
rect 418172 40174 418936 40202
rect 412836 40035 413120 40063
rect 413480 40038 413900 40066
rect 414308 40035 414680 40063
rect 415460 40035 415716 40063
rect 412836 27130 412864 40035
rect 412824 27124 412876 27130
rect 412824 27066 412876 27072
rect 414308 26234 414336 40035
rect 415688 38214 415716 40035
rect 415780 40035 416240 40063
rect 416792 40035 417020 40063
rect 417436 40035 417800 40063
rect 414664 38208 414716 38214
rect 414664 38150 414716 38156
rect 415676 38208 415728 38214
rect 415676 38150 415728 38156
rect 414032 26206 414336 26234
rect 412732 24336 412784 24342
rect 412732 24278 412784 24284
rect 414032 14482 414060 26206
rect 414020 14476 414072 14482
rect 414020 14418 414072 14424
rect 414676 13122 414704 38150
rect 415780 28354 415808 40035
rect 415768 28348 415820 28354
rect 415768 28290 415820 28296
rect 416792 17474 416820 40035
rect 417436 29850 417464 40035
rect 417424 29844 417476 29850
rect 417424 29786 417476 29792
rect 418172 22846 418200 40174
rect 418908 40066 418936 40174
rect 423692 40174 424180 40202
rect 418264 40035 418580 40063
rect 418908 40038 419360 40066
rect 419736 40035 420160 40063
rect 420940 40035 421052 40063
rect 418264 31278 418292 40035
rect 419736 35426 419764 40035
rect 420920 37868 420972 37874
rect 420920 37810 420972 37816
rect 419724 35420 419776 35426
rect 419724 35362 419776 35368
rect 418252 31272 418304 31278
rect 418252 31214 418304 31220
rect 419540 26988 419592 26994
rect 419540 26930 419592 26936
rect 418160 22840 418212 22846
rect 418160 22782 418212 22788
rect 416780 17468 416832 17474
rect 416780 17410 416832 17416
rect 419552 16574 419580 26930
rect 419552 16546 420224 16574
rect 417424 13320 417476 13326
rect 417424 13262 417476 13268
rect 414296 13116 414348 13122
rect 414296 13058 414348 13064
rect 414664 13116 414716 13122
rect 414664 13058 414716 13064
rect 414308 480 414336 13058
rect 415492 12028 415544 12034
rect 415492 11970 415544 11976
rect 415400 3664 415452 3670
rect 415400 3606 415452 3612
rect 415412 1850 415440 3606
rect 415504 3534 415532 11970
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 415412 1822 415532 1850
rect 415504 480 415532 1822
rect 416700 480 416728 3470
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 13262
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 419000 480 419028 3538
rect 420196 480 420224 16546
rect 420932 3602 420960 37810
rect 421024 25770 421052 40035
rect 421392 40035 421720 40063
rect 422480 40035 422800 40063
rect 421392 37874 421420 40035
rect 421380 37868 421432 37874
rect 421380 37810 421432 37816
rect 422772 36582 422800 40035
rect 422864 40035 423260 40063
rect 422760 36576 422812 36582
rect 422760 36518 422812 36524
rect 422864 26234 422892 40035
rect 422404 26206 422892 26234
rect 421012 25764 421064 25770
rect 421012 25706 421064 25712
rect 421012 13252 421064 13258
rect 421012 13194 421064 13200
rect 420920 3596 420972 3602
rect 420920 3538 420972 3544
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421024 354 421052 13194
rect 422404 3534 422432 26206
rect 423692 11626 423720 40174
rect 424152 40066 424180 40174
rect 428462 40080 428518 40089
rect 423784 40035 424040 40063
rect 424152 40038 424560 40066
rect 423784 12050 423812 40035
rect 428462 40015 428518 40024
rect 425704 38344 425756 38350
rect 425704 38286 425756 38292
rect 424968 13184 425020 13190
rect 424968 13126 425020 13132
rect 423784 12022 423996 12050
rect 423680 11620 423732 11626
rect 423680 11562 423732 11568
rect 423968 11506 423996 12022
rect 423692 11478 423996 11506
rect 423692 3754 423720 11478
rect 423772 11416 423824 11422
rect 423772 11358 423824 11364
rect 423600 3726 423720 3754
rect 423600 3670 423628 3726
rect 423588 3664 423640 3670
rect 423784 3618 423812 11358
rect 423864 10668 423916 10674
rect 423864 10610 423916 10616
rect 423588 3606 423640 3612
rect 423692 3590 423812 3618
rect 422392 3528 422444 3534
rect 422392 3470 422444 3476
rect 423692 3466 423720 3590
rect 423876 3482 423904 10610
rect 422576 3460 422628 3466
rect 422576 3402 422628 3408
rect 423680 3460 423732 3466
rect 423680 3402 423732 3408
rect 423784 3454 423904 3482
rect 422588 480 422616 3402
rect 423784 480 423812 3454
rect 424980 480 425008 13126
rect 425716 10674 425744 38286
rect 426440 29708 426492 29714
rect 426440 29650 426492 29656
rect 426452 16574 426480 29650
rect 427820 23112 427872 23118
rect 427820 23054 427872 23060
rect 426452 16546 426848 16574
rect 425704 10668 425756 10674
rect 425704 10610 425756 10616
rect 426164 3256 426216 3262
rect 426164 3198 426216 3204
rect 426176 480 426204 3198
rect 421350 354 421462 480
rect 421024 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 427832 6914 427860 23054
rect 428476 16574 428504 40015
rect 428568 20670 428596 48991
rect 428660 33114 428688 59327
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 447140 38276 447192 38282
rect 447140 38218 447192 38224
rect 436744 38208 436796 38214
rect 436744 38150 436796 38156
rect 434720 35556 434772 35562
rect 434720 35498 434772 35504
rect 428648 33108 428700 33114
rect 428648 33050 428700 33056
rect 428556 20664 428608 20670
rect 428556 20606 428608 20612
rect 432052 20120 432104 20126
rect 432052 20062 432104 20068
rect 430580 20052 430632 20058
rect 430580 19994 430632 20000
rect 430592 16574 430620 19994
rect 428476 16546 428596 16574
rect 430592 16546 430896 16574
rect 427832 6886 428504 6914
rect 428476 480 428504 6886
rect 428568 6866 428596 16546
rect 428556 6860 428608 6866
rect 428556 6802 428608 6808
rect 429660 3324 429712 3330
rect 429660 3266 429712 3272
rect 429672 480 429700 3266
rect 430868 480 430896 16546
rect 432064 480 432092 20062
rect 434732 16574 434760 35498
rect 434732 16546 435128 16574
rect 433984 10600 434036 10606
rect 433984 10542 434036 10548
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 10542
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 10606 436784 38150
rect 445760 32632 445812 32638
rect 445760 32574 445812 32580
rect 441620 31340 441672 31346
rect 441620 31282 441672 31288
rect 438860 17536 438912 17542
rect 438860 17478 438912 17484
rect 438872 16574 438900 17478
rect 441632 16574 441660 31282
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 436744 10600 436796 10606
rect 436744 10542 436796 10548
rect 437480 10532 437532 10538
rect 437480 10474 437532 10480
rect 436744 4140 436796 4146
rect 436744 4082 436796 4088
rect 436756 480 436784 4082
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 10474
rect 439148 480 439176 16546
rect 440332 10464 440384 10470
rect 440332 10406 440384 10412
rect 440240 4072 440292 4078
rect 440240 4014 440292 4020
rect 440252 2122 440280 4014
rect 440344 3398 440372 10406
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 2094 440372 2122
rect 440344 480 440372 2094
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 445024 10396 445076 10402
rect 445024 10338 445076 10344
rect 443828 4004 443880 4010
rect 443828 3946 443880 3952
rect 443840 480 443868 3946
rect 445036 480 445064 10338
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 32574
rect 447152 16574 447180 38218
rect 454040 38140 454092 38146
rect 454040 38082 454092 38088
rect 452660 27260 452712 27266
rect 452660 27202 452712 27208
rect 451280 25628 451332 25634
rect 451280 25570 451332 25576
rect 448520 18692 448572 18698
rect 448520 18634 448572 18640
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3210 448560 18634
rect 451292 16574 451320 25570
rect 452672 16574 452700 27202
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 16040 448664 16046
rect 448612 15982 448664 15988
rect 448624 3398 448652 15982
rect 450912 3936 450964 3942
rect 450912 3878 450964 3884
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 3878
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 38082
rect 460940 38072 460992 38078
rect 460940 38014 460992 38020
rect 458180 33924 458232 33930
rect 458180 33866 458232 33872
rect 456892 25832 456944 25838
rect 456892 25774 456944 25780
rect 455696 10328 455748 10334
rect 455696 10270 455748 10276
rect 455708 480 455736 10270
rect 456904 480 456932 25774
rect 458192 16574 458220 33866
rect 460952 16574 460980 38014
rect 467840 38004 467892 38010
rect 467840 37946 467892 37952
rect 466460 36780 466512 36786
rect 466460 36722 466512 36728
rect 465172 32496 465224 32502
rect 465172 32438 465224 32444
rect 463700 21684 463752 21690
rect 463700 21626 463752 21632
rect 462320 17400 462372 17406
rect 462320 17342 462372 17348
rect 458192 16546 459232 16574
rect 460952 16546 461624 16574
rect 458088 3868 458140 3874
rect 458088 3810 458140 3816
rect 458100 480 458128 3810
rect 459204 480 459232 16546
rect 459928 14748 459980 14754
rect 459928 14690 459980 14696
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 14690
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 17342
rect 463712 16574 463740 21626
rect 465184 16574 465212 32438
rect 466472 16574 466500 36722
rect 467852 16574 467880 37946
rect 474740 37936 474792 37942
rect 474740 37878 474792 37884
rect 469220 24200 469272 24206
rect 469220 24142 469272 24148
rect 469232 16574 469260 24142
rect 474752 16574 474780 37878
rect 538220 36712 538272 36718
rect 538220 36654 538272 36660
rect 534080 35352 534132 35358
rect 534080 35294 534132 35300
rect 483020 35284 483072 35290
rect 483020 35226 483072 35232
rect 476120 31204 476172 31210
rect 476120 31146 476172 31152
rect 476132 16574 476160 31146
rect 480260 17332 480312 17338
rect 480260 17274 480312 17280
rect 480272 16574 480300 17274
rect 483032 16574 483060 35226
rect 521660 33992 521712 33998
rect 521660 33934 521712 33940
rect 489920 33856 489972 33862
rect 489920 33798 489972 33804
rect 487160 18624 487212 18630
rect 487160 18566 487212 18572
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 480272 16546 480576 16574
rect 483032 16546 484072 16574
rect 463988 480 464016 16546
rect 465172 3800 465224 3806
rect 465172 3742 465224 3748
rect 465184 480 465212 3742
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 473452 16244 473504 16250
rect 473452 16186 473504 16192
rect 470600 14680 470652 14686
rect 470600 14622 470652 14628
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 14622
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473464 480 473492 16186
rect 474096 14612 474148 14618
rect 474096 14554 474148 14560
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 14554
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478144 14544 478196 14550
rect 478144 14486 478196 14492
rect 478156 480 478184 14486
rect 479338 3360 479394 3369
rect 479338 3295 479394 3304
rect 479352 480 479380 3295
rect 480548 480 480576 16546
rect 482836 9240 482888 9246
rect 482836 9182 482888 9188
rect 481732 6656 481784 6662
rect 481732 6598 481784 6604
rect 481744 480 481772 6598
rect 482848 480 482876 9182
rect 484044 480 484072 16546
rect 486424 9172 486476 9178
rect 486424 9114 486476 9120
rect 485228 6588 485280 6594
rect 485228 6530 485280 6536
rect 485240 480 485268 6530
rect 486436 480 486464 9114
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 18566
rect 489932 16574 489960 33798
rect 494060 31136 494112 31142
rect 494060 31078 494112 31084
rect 494072 16574 494100 31078
rect 506480 29912 506532 29918
rect 506480 29854 506532 29860
rect 500960 29640 501012 29646
rect 500960 29582 501012 29588
rect 499580 28484 499632 28490
rect 499580 28426 499632 28432
rect 498200 21412 498252 21418
rect 498200 21354 498252 21360
rect 489932 16546 490696 16574
rect 494072 16546 494744 16574
rect 489920 9104 489972 9110
rect 489920 9046 489972 9052
rect 488816 6520 488868 6526
rect 488816 6462 488868 6468
rect 488828 480 488856 6462
rect 489932 480 489960 9046
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 493508 9036 493560 9042
rect 493508 8978 493560 8984
rect 492312 6452 492364 6458
rect 492312 6394 492364 6400
rect 492324 480 492352 6394
rect 493520 480 493548 8978
rect 494716 480 494744 16546
rect 497096 8968 497148 8974
rect 497096 8910 497148 8916
rect 495900 6384 495952 6390
rect 495900 6326 495952 6332
rect 495912 480 495940 6326
rect 497108 480 497136 8910
rect 498212 480 498240 21354
rect 499592 16574 499620 28426
rect 500972 16574 501000 29582
rect 505100 22772 505152 22778
rect 505100 22714 505152 22720
rect 505112 16574 505140 22714
rect 506492 16574 506520 29854
rect 513380 28416 513432 28422
rect 513380 28358 513432 28364
rect 507860 28280 507912 28286
rect 507860 28222 507912 28228
rect 507872 16574 507900 28222
rect 512000 26920 512052 26926
rect 512000 26862 512052 26868
rect 509240 21548 509292 21554
rect 509240 21490 509292 21496
rect 509252 16574 509280 21490
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 505112 16546 505416 16574
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 499396 6316 499448 6322
rect 499396 6258 499448 6264
rect 499408 480 499436 6258
rect 500604 480 500632 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 503720 13524 503772 13530
rect 503720 13466 503772 13472
rect 502984 6248 503036 6254
rect 502984 6190 503036 6196
rect 502996 480 503024 6190
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 13466
rect 505388 480 505416 16546
rect 506480 6180 506532 6186
rect 506480 6122 506532 6128
rect 506492 480 506520 6122
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 11892 511316 11898
rect 511264 11834 511316 11840
rect 511276 480 511304 11834
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 26862
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 28358
rect 520280 27056 520332 27062
rect 520280 26998 520332 27004
rect 514760 22976 514812 22982
rect 514760 22918 514812 22924
rect 514772 480 514800 22918
rect 516140 22908 516192 22914
rect 516140 22850 516192 22856
rect 516152 16574 516180 22850
rect 517520 18828 517572 18834
rect 517520 18770 517572 18776
rect 517532 16574 517560 18770
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 515956 5228 516008 5234
rect 515956 5170 516008 5176
rect 515968 480 515996 5170
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 5160 519596 5166
rect 519544 5102 519596 5108
rect 519556 480 519584 5102
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 26998
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 33934
rect 523040 29776 523092 29782
rect 523040 29718 523092 29724
rect 523052 3398 523080 29718
rect 523132 24132 523184 24138
rect 523132 24074 523184 24080
rect 523040 3392 523092 3398
rect 523040 3334 523092 3340
rect 523144 3210 523172 24074
rect 528560 21480 528612 21486
rect 528560 21422 528612 21428
rect 524420 20188 524472 20194
rect 524420 20130 524472 20136
rect 524432 16574 524460 20130
rect 527180 18760 527232 18766
rect 527180 18702 527232 18708
rect 527192 16574 527220 18702
rect 524432 16546 525472 16574
rect 527192 16546 527864 16574
rect 523868 3392 523920 3398
rect 523868 3334 523920 3340
rect 523052 3182 523172 3210
rect 523052 480 523080 3182
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3334
rect 525444 480 525472 16546
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526640 480 526668 5034
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 21422
rect 534092 16574 534120 35294
rect 534092 16546 534488 16574
rect 531320 11824 531372 11830
rect 531320 11766 531372 11772
rect 530124 5024 530176 5030
rect 530124 4966 530176 4972
rect 530136 480 530164 4966
rect 531332 480 531360 11766
rect 532056 10668 532108 10674
rect 532056 10610 532108 10616
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 10610
rect 533712 4956 533764 4962
rect 533712 4898 533764 4904
rect 533724 480 533752 4898
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536104 13388 536156 13394
rect 536104 13330 536156 13336
rect 536116 480 536144 13330
rect 537208 4888 537260 4894
rect 537208 4830 537260 4836
rect 537220 480 537248 4830
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 36654
rect 557540 36644 557592 36650
rect 557540 36586 557592 36592
rect 554780 32428 554832 32434
rect 554780 32370 554832 32376
rect 553400 28348 553452 28354
rect 553400 28290 553452 28296
rect 539600 27124 539652 27130
rect 539600 27066 539652 27072
rect 539612 480 539640 27066
rect 547880 25696 547932 25702
rect 547880 25638 547932 25644
rect 543740 25560 543792 25566
rect 543740 25502 543792 25508
rect 542360 24336 542412 24342
rect 542360 24278 542412 24284
rect 542372 16574 542400 24278
rect 543752 16574 543780 25502
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 541992 8016 542044 8022
rect 541992 7958 542044 7964
rect 540796 4820 540848 4826
rect 540796 4762 540848 4768
rect 540808 480 540836 4762
rect 542004 480 542032 7958
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 15904 545540 15910
rect 545488 15846 545540 15852
rect 545500 480 545528 15846
rect 546500 14476 546552 14482
rect 546500 14418 546552 14424
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 14418
rect 547892 3398 547920 25638
rect 550640 19984 550692 19990
rect 550640 19926 550692 19932
rect 550652 16574 550680 19926
rect 553412 16574 553440 28290
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 547972 15972 548024 15978
rect 547972 15914 548024 15920
rect 547880 3392 547932 3398
rect 547880 3334 547932 3340
rect 547984 3210 548012 15914
rect 550272 10600 550324 10606
rect 550272 10542 550324 10548
rect 548708 3392 548760 3398
rect 548708 3334 548760 3340
rect 547892 3182 548012 3210
rect 547892 480 547920 3182
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3334
rect 550284 480 550312 10542
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 7948 552716 7954
rect 552664 7890 552716 7896
rect 552676 480 552704 7890
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 32370
rect 556160 17468 556212 17474
rect 556160 17410 556212 17416
rect 556172 16574 556200 17410
rect 557552 16574 557580 36586
rect 579620 36576 579672 36582
rect 579620 36518 579672 36524
rect 571340 35420 571392 35426
rect 571340 35362 571392 35368
rect 564440 35216 564492 35222
rect 564440 35158 564492 35164
rect 560300 29844 560352 29850
rect 560300 29786 560352 29792
rect 560312 16574 560340 29786
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 556160 7880 556212 7886
rect 556160 7822 556212 7828
rect 556172 480 556200 7822
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 559748 7812 559800 7818
rect 559748 7754 559800 7760
rect 559760 480 559788 7754
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 562048 11756 562100 11762
rect 562048 11698 562100 11704
rect 562060 480 562088 11698
rect 563244 7744 563296 7750
rect 563244 7686 563296 7692
rect 563256 480 563284 7686
rect 564452 3398 564480 35158
rect 564532 31272 564584 31278
rect 564532 31214 564584 31220
rect 564440 3392 564492 3398
rect 564440 3334 564492 3340
rect 564544 3210 564572 31214
rect 565820 24268 565872 24274
rect 565820 24210 565872 24216
rect 565832 16574 565860 24210
rect 567200 22840 567252 22846
rect 567200 22782 567252 22788
rect 567212 16574 567240 22782
rect 568580 17264 568632 17270
rect 568580 17206 568632 17212
rect 568592 16574 568620 17206
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 565268 3392 565320 3398
rect 565268 3334 565320 3340
rect 564452 3182 564572 3210
rect 564452 480 564480 3182
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565280 354 565308 3334
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570328 7676 570380 7682
rect 570328 7618 570380 7624
rect 570340 480 570368 7618
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 35362
rect 572720 33788 572772 33794
rect 572720 33730 572772 33736
rect 572732 480 572760 33730
rect 575480 31068 575532 31074
rect 575480 31010 575532 31016
rect 574100 25764 574152 25770
rect 574100 25706 574152 25712
rect 574112 16574 574140 25706
rect 575492 16574 575520 31010
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 573916 7608 573968 7614
rect 573916 7550 573968 7556
rect 573928 480 573956 7550
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576952 13116 577004 13122
rect 576952 13058 577004 13064
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 13058
rect 578608 3596 578660 3602
rect 578608 3538 578660 3544
rect 578620 480 578648 3538
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579632 354 579660 36518
rect 579894 33144 579950 33153
rect 579894 33079 579896 33088
rect 579948 33079 579950 33088
rect 579896 33050 579948 33056
rect 579896 20664 579948 20670
rect 579896 20606 579948 20612
rect 579908 19825 579936 20606
rect 579894 19816 579950 19825
rect 579894 19751 579950 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 582196 3664 582248 3670
rect 582196 3606 582248 3612
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 582208 480 582236 3606
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3514 684256 3570 684312
rect 3422 671200 3478 671256
rect 2870 645088 2926 645144
rect 3330 606056 3386 606112
rect 3330 593000 3386 593056
rect 3330 579944 3386 580000
rect 3146 553832 3202 553888
rect 3054 540776 3110 540832
rect 2962 527856 3018 527912
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3422 514800 3478 514856
rect 3146 488688 3202 488744
rect 3330 436600 3386 436656
rect 3330 423544 3386 423600
rect 3606 566888 3662 566944
rect 3514 475632 3570 475688
rect 3514 462576 3570 462632
rect 3422 410488 3478 410544
rect 3330 384376 3386 384432
rect 3146 371340 3202 371376
rect 3146 371320 3148 371340
rect 3148 371320 3200 371340
rect 3200 371320 3202 371340
rect 3698 501744 3754 501800
rect 3790 449520 3846 449576
rect 3606 397432 3662 397488
rect 3514 358400 3570 358456
rect 2778 332288 2834 332344
rect 3422 319232 3478 319288
rect 3698 345344 3754 345400
rect 3606 306176 3662 306232
rect 3514 293120 3570 293176
rect 3422 267144 3478 267200
rect 3698 280064 3754 280120
rect 3606 254088 3662 254144
rect 3514 241032 3570 241088
rect 3422 227976 3478 228032
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 37830 544584 37886 544640
rect 37554 536152 37610 536208
rect 37830 526632 37886 526688
rect 37554 507456 37610 507512
rect 579618 630808 579674 630864
rect 428462 535336 428518 535392
rect 38014 517112 38070 517168
rect 37922 498072 37978 498128
rect 37830 488452 37832 488472
rect 37832 488452 37884 488472
rect 37884 488452 37886 488472
rect 37830 488416 37886 488452
rect 36542 478352 36598 478408
rect 37922 468832 37978 468888
rect 37462 459312 37518 459368
rect 37922 449828 37924 449848
rect 37924 449828 37976 449848
rect 37976 449828 37978 449848
rect 37922 449792 37978 449828
rect 37830 440816 37886 440872
rect 37830 431296 37886 431352
rect 37922 421776 37978 421832
rect 580170 577632 580226 577688
rect 428554 496712 428610 496768
rect 428554 487092 428556 487112
rect 428556 487092 428608 487112
rect 428608 487092 428610 487112
rect 428554 487056 428610 487092
rect 428554 477436 428556 477456
rect 428556 477436 428608 477456
rect 428608 477436 428610 477456
rect 428554 477400 428610 477436
rect 428462 419464 428518 419520
rect 37646 412256 37702 412312
rect 37554 402464 37610 402520
rect 428462 399880 428518 399936
rect 37738 393080 37794 393136
rect 428462 390088 428518 390144
rect 37462 383596 37464 383616
rect 37464 383596 37516 383616
rect 37516 383596 37518 383616
rect 37462 383560 37518 383596
rect 580170 551112 580226 551168
rect 428738 544856 428794 544912
rect 428738 525716 428740 525736
rect 428740 525716 428792 525736
rect 428792 525716 428794 525736
rect 428738 525680 428794 525716
rect 428738 516060 428740 516080
rect 428740 516060 428792 516080
rect 428792 516060 428794 516080
rect 428738 516024 428794 516060
rect 428738 506404 428740 506424
rect 428740 506404 428792 506424
rect 428792 506404 428794 506424
rect 428738 506368 428794 506404
rect 428738 467780 428740 467800
rect 428740 467780 428792 467800
rect 428792 467780 428794 467800
rect 428738 467744 428794 467780
rect 428646 458088 428702 458144
rect 429106 448160 429162 448216
rect 580354 670656 580410 670712
rect 580262 537784 580318 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 579986 471416 580042 471472
rect 428646 438640 428702 438696
rect 580078 431568 580134 431624
rect 428646 428984 428702 429040
rect 580446 657328 580502 657384
rect 580538 644000 580594 644056
rect 580354 511264 580410 511320
rect 428554 380568 428610 380624
rect 37922 373940 37924 373960
rect 37924 373940 37976 373960
rect 37976 373940 37978 373960
rect 37922 373904 37978 373940
rect 37462 364112 37518 364168
rect 37554 354456 37610 354512
rect 37646 344972 37648 344992
rect 37648 344972 37700 344992
rect 37700 344972 37702 344992
rect 37646 344936 37702 344972
rect 37830 335960 37886 336016
rect 37554 326440 37610 326496
rect 37922 316920 37978 316976
rect 37370 307264 37426 307320
rect 428554 361120 428610 361176
rect 580170 418240 580226 418296
rect 428646 351328 428702 351384
rect 580630 617480 580686 617536
rect 580446 497936 580502 497992
rect 428830 409400 428886 409456
rect 580262 404912 580318 404968
rect 428830 370640 428886 370696
rect 579802 365064 579858 365120
rect 428738 341672 428794 341728
rect 580722 604152 580778 604208
rect 580538 484608 580594 484664
rect 580354 391720 580410 391776
rect 428554 332016 428610 332072
rect 579618 325216 579674 325272
rect 428462 302776 428518 302832
rect 37554 297608 37610 297664
rect 428462 292476 428464 292496
rect 428464 292476 428516 292496
rect 428516 292476 428518 292496
rect 428462 292440 428518 292476
rect 37738 288224 37794 288280
rect 37738 278432 37794 278488
rect 580814 590960 580870 591016
rect 580906 564304 580962 564360
rect 580630 458088 580686 458144
rect 580446 378392 580502 378448
rect 428830 322224 428886 322280
rect 580722 444760 580778 444816
rect 580538 351872 580594 351928
rect 428738 312568 428794 312624
rect 580170 312024 580226 312080
rect 428554 273128 428610 273184
rect 37922 268912 37978 268968
rect 37370 258032 37426 258088
rect 37922 249600 37978 249656
rect 37370 240100 37426 240136
rect 37370 240080 37372 240100
rect 37372 240080 37424 240100
rect 37424 240080 37426 240100
rect 580262 298696 580318 298752
rect 429014 282820 429016 282840
rect 429016 282820 429068 282840
rect 429068 282820 429070 282840
rect 429014 282784 429070 282820
rect 579618 272176 579674 272232
rect 428646 263472 428702 263528
rect 579618 258848 579674 258904
rect 428462 234504 428518 234560
rect 37646 230560 37702 230616
rect 37738 221584 37794 221640
rect 3606 214920 3662 214976
rect 3514 201864 3570 201920
rect 3422 188808 3478 188864
rect 37830 212064 37886 212120
rect 580630 338544 580686 338600
rect 580354 285368 580410 285424
rect 428922 253852 428924 253872
rect 428924 253852 428976 253872
rect 428976 253852 428978 253872
rect 428922 253816 428978 253852
rect 579802 245520 579858 245576
rect 428646 244196 428648 244216
rect 428648 244196 428700 244216
rect 428700 244196 428702 244216
rect 428646 244160 428702 244196
rect 428554 224848 428610 224904
rect 428462 205536 428518 205592
rect 37738 202544 37794 202600
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 428646 215192 428702 215248
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 428554 195880 428610 195936
rect 37738 192888 37794 192944
rect 37922 183368 37978 183424
rect 580170 192480 580226 192536
rect 428646 186224 428702 186280
rect 580170 179152 580226 179208
rect 428462 176568 428518 176624
rect 3514 175888 3570 175944
rect 37738 173576 37794 173632
rect 428554 166776 428610 166832
rect 580170 165824 580226 165880
rect 37922 164056 37978 164112
rect 3422 162832 3478 162888
rect 428462 157120 428518 157176
rect 37646 154264 37702 154320
rect 579986 152632 580042 152688
rect 3330 149776 3386 149832
rect 429106 147328 429162 147384
rect 37922 144744 37978 144800
rect 580170 139304 580226 139360
rect 428830 137536 428886 137592
rect 3422 136720 3478 136776
rect 37554 135768 37610 135824
rect 428922 127064 428978 127120
rect 580170 125976 580226 126032
rect 37738 125704 37794 125760
rect 3422 123664 3478 123720
rect 428462 117272 428518 117328
rect 37922 115912 37978 115968
rect 579802 112784 579858 112840
rect 3422 110608 3478 110664
rect 428462 107616 428518 107672
rect 37922 106256 37978 106312
rect 580170 99456 580226 99512
rect 428554 97960 428610 98016
rect 3422 97552 3478 97608
rect 38014 96600 38070 96656
rect 37922 86944 37978 87000
rect 3146 84632 3202 84688
rect 428462 88304 428518 88360
rect 38014 77424 38070 77480
rect 3422 71576 3478 71632
rect 37922 67904 37978 67960
rect 3054 58520 3110 58576
rect 580170 86128 580226 86184
rect 428554 78648 428610 78704
rect 428462 69128 428518 69184
rect 38106 58384 38162 58440
rect 38014 49272 38070 49328
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 37922 40160 37978 40216
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 428646 59336 428702 59392
rect 428554 49000 428610 49056
rect 120262 3304 120318 3360
rect 305550 3304 305606 3360
rect 361578 3304 361634 3360
rect 398838 3304 398894 3360
rect 428462 40024 428518 40080
rect 580170 46280 580226 46336
rect 479338 3304 479394 3360
rect 579894 33108 579950 33144
rect 579894 33088 579896 33108
rect 579896 33088 579948 33108
rect 579948 33088 579950 33108
rect 579894 19760 579950 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580349 670714 580415 670717
rect 583520 670714 584960 670804
rect 580349 670712 584960 670714
rect 580349 670656 580354 670712
rect 580410 670656 584960 670712
rect 580349 670654 584960 670656
rect 580349 670651 580415 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 580441 657386 580507 657389
rect 583520 657386 584960 657476
rect 580441 657384 584960 657386
rect 580441 657328 580446 657384
rect 580502 657328 584960 657384
rect 580441 657326 584960 657328
rect 580441 657323 580507 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 2865 645146 2931 645149
rect -960 645144 2931 645146
rect -960 645088 2870 645144
rect 2926 645088 2931 645144
rect -960 645086 2931 645088
rect -960 644996 480 645086
rect 2865 645083 2931 645086
rect 580533 644058 580599 644061
rect 583520 644058 584960 644148
rect 580533 644056 584960 644058
rect 580533 644000 580538 644056
rect 580594 644000 584960 644056
rect 580533 643998 584960 644000
rect 580533 643995 580599 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 579613 630866 579679 630869
rect 583520 630866 584960 630956
rect 579613 630864 584960 630866
rect 579613 630808 579618 630864
rect 579674 630808 584960 630864
rect 579613 630806 584960 630808
rect 579613 630803 579679 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580625 617538 580691 617541
rect 583520 617538 584960 617628
rect 580625 617536 584960 617538
rect 580625 617480 580630 617536
rect 580686 617480 584960 617536
rect 580625 617478 584960 617480
rect 580625 617475 580691 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 580717 604210 580783 604213
rect 583520 604210 584960 604300
rect 580717 604208 584960 604210
rect 580717 604152 580722 604208
rect 580778 604152 584960 604208
rect 580717 604150 584960 604152
rect 580717 604147 580783 604150
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3325 593058 3391 593061
rect -960 593056 3391 593058
rect -960 593000 3330 593056
rect 3386 593000 3391 593056
rect -960 592998 3391 593000
rect -960 592908 480 592998
rect 3325 592995 3391 592998
rect 580809 591018 580875 591021
rect 583520 591018 584960 591108
rect 580809 591016 584960 591018
rect 580809 590960 580814 591016
rect 580870 590960 584960 591016
rect 580809 590958 584960 590960
rect 580809 590955 580875 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 580901 564362 580967 564365
rect 583520 564362 584960 564452
rect 580901 564360 584960 564362
rect 580901 564304 580906 564360
rect 580962 564304 584960 564360
rect 580901 564302 584960 564304
rect 580901 564299 580967 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 580165 551170 580231 551173
rect 583520 551170 584960 551260
rect 580165 551168 584960 551170
rect 580165 551112 580170 551168
rect 580226 551112 584960 551168
rect 580165 551110 584960 551112
rect 580165 551107 580231 551110
rect 583520 551020 584960 551110
rect 428733 544914 428799 544917
rect 425194 544912 428799 544914
rect 425194 544856 428738 544912
rect 428794 544856 428799 544912
rect 425194 544854 428799 544856
rect 425194 544710 425254 544854
rect 428733 544851 428799 544854
rect 37825 544642 37891 544645
rect 37825 544640 39498 544642
rect 37825 544584 37830 544640
rect 37886 544625 39498 544640
rect 37886 544584 40020 544625
rect 37825 544582 40020 544584
rect 37825 544579 37891 544582
rect 39438 544565 40020 544582
rect -960 540834 480 540924
rect 3049 540834 3115 540837
rect -960 540832 3115 540834
rect -960 540776 3054 540832
rect 3110 540776 3115 540832
rect -960 540774 3115 540776
rect -960 540684 480 540774
rect 3049 540771 3115 540774
rect 580257 537842 580323 537845
rect 583520 537842 584960 537932
rect 580257 537840 584960 537842
rect 580257 537784 580262 537840
rect 580318 537784 584960 537840
rect 580257 537782 584960 537784
rect 580257 537779 580323 537782
rect 583520 537692 584960 537782
rect 37549 536210 37615 536213
rect 37549 536208 40110 536210
rect 37549 536152 37554 536208
rect 37610 536152 40110 536208
rect 37549 536150 40110 536152
rect 37549 536147 37615 536150
rect 40050 535571 40110 536150
rect 425194 535394 425254 535398
rect 428457 535394 428523 535397
rect 425194 535392 428523 535394
rect 425194 535336 428462 535392
rect 428518 535336 428523 535392
rect 425194 535334 428523 535336
rect 428457 535331 428523 535334
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 37825 526690 37891 526693
rect 37825 526688 40110 526690
rect 37825 526632 37830 526688
rect 37886 526632 40110 526688
rect 37825 526630 40110 526632
rect 37825 526627 37891 526630
rect 40050 526067 40110 526630
rect 428733 525738 428799 525741
rect 425194 525736 428799 525738
rect 425194 525680 428738 525736
rect 428794 525680 428799 525736
rect 425194 525678 428799 525680
rect 428733 525675 428799 525678
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 38009 517170 38075 517173
rect 38009 517168 40110 517170
rect 38009 517112 38014 517168
rect 38070 517112 40110 517168
rect 38009 517110 40110 517112
rect 38009 517107 38075 517110
rect 40050 516525 40110 517110
rect 428733 516082 428799 516085
rect 425838 516080 428799 516082
rect 425838 516024 428738 516080
rect 428794 516024 428799 516080
rect 425838 516022 428799 516024
rect 425838 516017 425898 516022
rect 428733 516019 428799 516022
rect 425224 515957 425898 516017
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580349 511322 580415 511325
rect 583520 511322 584960 511412
rect 580349 511320 584960 511322
rect 580349 511264 580354 511320
rect 580410 511264 584960 511320
rect 580349 511262 584960 511264
rect 580349 511259 580415 511262
rect 583520 511172 584960 511262
rect 37549 507514 37615 507517
rect 37549 507512 40110 507514
rect 37549 507456 37554 507512
rect 37610 507456 40110 507512
rect 37549 507454 40110 507456
rect 37549 507451 37615 507454
rect 40050 506963 40110 507454
rect 428733 506426 428799 506429
rect 425194 506424 428799 506426
rect 425194 506368 428738 506424
rect 428794 506368 428799 506424
rect 425194 506366 428799 506368
rect 425194 506253 425254 506366
rect 428733 506363 428799 506366
rect -960 501802 480 501892
rect 3693 501802 3759 501805
rect -960 501800 3759 501802
rect -960 501744 3698 501800
rect 3754 501744 3759 501800
rect -960 501742 3759 501744
rect -960 501652 480 501742
rect 3693 501739 3759 501742
rect 37917 498130 37983 498133
rect 37917 498128 40110 498130
rect 37917 498072 37922 498128
rect 37978 498072 40110 498128
rect 37917 498070 40110 498072
rect 37917 498067 37983 498070
rect 40050 497459 40110 498070
rect 580441 497994 580507 497997
rect 583520 497994 584960 498084
rect 580441 497992 584960 497994
rect 580441 497936 580446 497992
rect 580502 497936 584960 497992
rect 580441 497934 584960 497936
rect 580441 497931 580507 497934
rect 583520 497844 584960 497934
rect 428549 496770 428615 496773
rect 425194 496768 428615 496770
rect 425194 496712 428554 496768
rect 428610 496712 428615 496768
rect 425194 496710 428615 496712
rect 425194 496518 425254 496710
rect 428549 496707 428615 496710
rect -960 488746 480 488836
rect 3141 488746 3207 488749
rect -960 488744 3207 488746
rect -960 488688 3146 488744
rect 3202 488688 3207 488744
rect -960 488686 3207 488688
rect -960 488596 480 488686
rect 3141 488683 3207 488686
rect 37825 488474 37891 488477
rect 37825 488472 40110 488474
rect 37825 488416 37830 488472
rect 37886 488416 40110 488472
rect 37825 488414 40110 488416
rect 37825 488411 37891 488414
rect 40050 487917 40110 488414
rect 428549 487114 428615 487117
rect 425194 487112 428615 487114
rect 425194 487056 428554 487112
rect 428610 487056 428615 487112
rect 425194 487054 428615 487056
rect 425194 486803 425254 487054
rect 428549 487051 428615 487054
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect 36537 478410 36603 478413
rect 39438 478410 40020 478424
rect 36537 478408 40020 478410
rect 36537 478352 36542 478408
rect 36598 478364 40020 478408
rect 36598 478352 39498 478364
rect 36537 478350 39498 478352
rect 36537 478347 36603 478350
rect 428549 477458 428615 477461
rect 425194 477456 428615 477458
rect 425194 477400 428554 477456
rect 428610 477400 428615 477456
rect 425194 477398 428615 477400
rect 425194 477107 425254 477398
rect 428549 477395 428615 477398
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 37917 468890 37983 468893
rect 37917 468888 39498 468890
rect 37917 468832 37922 468888
rect 37978 468881 39498 468888
rect 37978 468832 40020 468881
rect 37917 468830 40020 468832
rect 37917 468827 37983 468830
rect 39438 468821 40020 468830
rect 428733 467802 428799 467805
rect 425186 467800 428799 467802
rect 425186 467744 428738 467800
rect 428794 467744 428799 467800
rect 425186 467742 428799 467744
rect 425186 467392 425246 467742
rect 428733 467739 428799 467742
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 37457 459370 37523 459373
rect 37457 459368 39498 459370
rect 37457 459312 37462 459368
rect 37518 459358 39498 459368
rect 37518 459312 40020 459358
rect 37457 459310 40020 459312
rect 37457 459307 37523 459310
rect 39438 459298 40020 459310
rect 428641 458146 428707 458149
rect 425194 458144 428707 458146
rect 425194 458088 428646 458144
rect 428702 458088 428707 458144
rect 425194 458086 428707 458088
rect 425194 457658 425254 458086
rect 428641 458083 428707 458086
rect 580625 458146 580691 458149
rect 583520 458146 584960 458236
rect 580625 458144 584960 458146
rect 580625 458088 580630 458144
rect 580686 458088 584960 458144
rect 580625 458086 584960 458088
rect 580625 458083 580691 458086
rect 583520 457996 584960 458086
rect 37917 449850 37983 449853
rect 37917 449848 40110 449850
rect 37917 449792 37922 449848
rect 37978 449792 40110 449848
rect 37917 449790 40110 449792
rect 37917 449787 37983 449790
rect 40050 449766 40110 449790
rect -960 449578 480 449668
rect 3785 449578 3851 449581
rect -960 449576 3851 449578
rect -960 449520 3790 449576
rect 3846 449520 3851 449576
rect -960 449518 3851 449520
rect -960 449428 480 449518
rect 3785 449515 3851 449518
rect 429101 448218 429167 448221
rect 425194 448216 429167 448218
rect 425194 448160 429106 448216
rect 429162 448160 429167 448216
rect 425194 448158 429167 448160
rect 425194 447962 425254 448158
rect 429101 448155 429167 448158
rect 580717 444818 580783 444821
rect 583520 444818 584960 444908
rect 580717 444816 584960 444818
rect 580717 444760 580722 444816
rect 580778 444760 584960 444816
rect 580717 444758 584960 444760
rect 580717 444755 580783 444758
rect 583520 444668 584960 444758
rect 37825 440874 37891 440877
rect 37825 440872 40110 440874
rect 37825 440816 37830 440872
rect 37886 440816 40110 440872
rect 37825 440814 40110 440816
rect 37825 440811 37891 440814
rect 40050 440262 40110 440814
rect 428641 438698 428707 438701
rect 425194 438696 428707 438698
rect 425194 438640 428646 438696
rect 428702 438640 428707 438696
rect 425194 438638 428707 438640
rect 425194 438246 425254 438638
rect 428641 438635 428707 438638
rect -960 436658 480 436748
rect 3325 436658 3391 436661
rect -960 436656 3391 436658
rect -960 436600 3330 436656
rect 3386 436600 3391 436656
rect -960 436598 3391 436600
rect -960 436508 480 436598
rect 3325 436595 3391 436598
rect 580073 431626 580139 431629
rect 583520 431626 584960 431716
rect 580073 431624 584960 431626
rect 580073 431568 580078 431624
rect 580134 431568 584960 431624
rect 580073 431566 584960 431568
rect 580073 431563 580139 431566
rect 583520 431476 584960 431566
rect 37825 431354 37891 431357
rect 37825 431352 40110 431354
rect 37825 431296 37830 431352
rect 37886 431296 40110 431352
rect 37825 431294 40110 431296
rect 37825 431291 37891 431294
rect 40050 430720 40110 431294
rect 428641 429042 428707 429045
rect 425194 429040 428707 429042
rect 425194 428984 428646 429040
rect 428702 428984 428707 429040
rect 425194 428982 428707 428984
rect 425194 428531 425254 428982
rect 428641 428979 428707 428982
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 37917 421834 37983 421837
rect 37917 421832 40110 421834
rect 37917 421776 37922 421832
rect 37978 421776 40110 421832
rect 37917 421774 40110 421776
rect 37917 421771 37983 421774
rect 40050 421197 40110 421774
rect 428457 419522 428523 419525
rect 425194 419520 428523 419522
rect 425194 419464 428462 419520
rect 428518 419464 428523 419520
rect 425194 419462 428523 419464
rect 425194 418854 425254 419462
rect 428457 419459 428523 419462
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 37641 412314 37707 412317
rect 37641 412312 40110 412314
rect 37641 412256 37646 412312
rect 37702 412256 40110 412312
rect 37641 412254 40110 412256
rect 37641 412251 37707 412254
rect 40050 411674 40110 412254
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 428825 409458 428891 409461
rect 425194 409456 428891 409458
rect 425194 409400 428830 409456
rect 428886 409400 428891 409456
rect 425194 409398 428891 409400
rect 425194 409101 425254 409398
rect 428825 409395 428891 409398
rect 580257 404970 580323 404973
rect 583520 404970 584960 405060
rect 580257 404968 584960 404970
rect 580257 404912 580262 404968
rect 580318 404912 584960 404968
rect 580257 404910 584960 404912
rect 580257 404907 580323 404910
rect 583520 404820 584960 404910
rect 37549 402522 37615 402525
rect 37549 402520 40110 402522
rect 37549 402464 37554 402520
rect 37610 402464 40110 402520
rect 37549 402462 40110 402464
rect 37549 402459 37615 402462
rect 40050 402131 40110 402462
rect 428457 399938 428523 399941
rect 425194 399936 428523 399938
rect 425194 399880 428462 399936
rect 428518 399880 428523 399936
rect 425194 399878 428523 399880
rect 425194 399386 425254 399878
rect 428457 399875 428523 399878
rect -960 397490 480 397580
rect 3601 397490 3667 397493
rect -960 397488 3667 397490
rect -960 397432 3606 397488
rect 3662 397432 3667 397488
rect -960 397430 3667 397432
rect -960 397340 480 397430
rect 3601 397427 3667 397430
rect 37733 393138 37799 393141
rect 37733 393136 40110 393138
rect 37733 393080 37738 393136
rect 37794 393080 40110 393136
rect 37733 393078 40110 393080
rect 37733 393075 37799 393078
rect 40050 392608 40110 393078
rect 580349 391778 580415 391781
rect 583520 391778 584960 391868
rect 580349 391776 584960 391778
rect 580349 391720 580354 391776
rect 580410 391720 584960 391776
rect 580349 391718 584960 391720
rect 580349 391715 580415 391718
rect 583520 391628 584960 391718
rect 428457 390146 428523 390149
rect 425194 390144 428523 390146
rect 425194 390088 428462 390144
rect 428518 390088 428523 390144
rect 425194 390086 428523 390088
rect 425194 389670 425254 390086
rect 428457 390083 428523 390086
rect -960 384434 480 384524
rect 3325 384434 3391 384437
rect -960 384432 3391 384434
rect -960 384376 3330 384432
rect 3386 384376 3391 384432
rect -960 384374 3391 384376
rect -960 384284 480 384374
rect 3325 384371 3391 384374
rect 37457 383618 37523 383621
rect 37457 383616 40110 383618
rect 37457 383560 37462 383616
rect 37518 383560 40110 383616
rect 37457 383558 40110 383560
rect 37457 383555 37523 383558
rect 40050 383066 40110 383558
rect 428549 380626 428615 380629
rect 425194 380624 428615 380626
rect 425194 380568 428554 380624
rect 428610 380568 428615 380624
rect 425194 380566 428615 380568
rect 425194 379974 425254 380566
rect 428549 380563 428615 380566
rect 580441 378450 580507 378453
rect 583520 378450 584960 378540
rect 580441 378448 584960 378450
rect 580441 378392 580446 378448
rect 580502 378392 584960 378448
rect 580441 378390 584960 378392
rect 580441 378387 580507 378390
rect 583520 378300 584960 378390
rect 37917 373962 37983 373965
rect 37917 373960 40110 373962
rect 37917 373904 37922 373960
rect 37978 373904 40110 373960
rect 37917 373902 40110 373904
rect 37917 373899 37983 373902
rect 40050 373562 40110 373902
rect -960 371378 480 371468
rect 3141 371378 3207 371381
rect -960 371376 3207 371378
rect -960 371320 3146 371376
rect 3202 371320 3207 371376
rect -960 371318 3207 371320
rect -960 371228 480 371318
rect 3141 371315 3207 371318
rect 428825 370698 428891 370701
rect 425194 370696 428891 370698
rect 425194 370640 428830 370696
rect 428886 370640 428891 370696
rect 425194 370638 428891 370640
rect 425194 370240 425254 370638
rect 428825 370635 428891 370638
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect 37457 364170 37523 364173
rect 37457 364168 40110 364170
rect 37457 364112 37462 364168
rect 37518 364112 40110 364168
rect 37457 364110 40110 364112
rect 37457 364107 37523 364110
rect 40050 364019 40110 364110
rect 428549 361178 428615 361181
rect 425194 361176 428615 361178
rect 425194 361120 428554 361176
rect 428610 361120 428615 361176
rect 425194 361118 428615 361120
rect 425194 360506 425254 361118
rect 428549 361115 428615 361118
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 37549 354514 37615 354517
rect 39438 354514 40020 354526
rect 37549 354512 40020 354514
rect 37549 354456 37554 354512
rect 37610 354466 40020 354512
rect 37610 354456 39498 354466
rect 37549 354454 39498 354456
rect 37549 354451 37615 354454
rect 580533 351930 580599 351933
rect 583520 351930 584960 352020
rect 580533 351928 584960 351930
rect 580533 351872 580538 351928
rect 580594 351872 584960 351928
rect 580533 351870 584960 351872
rect 580533 351867 580599 351870
rect 583520 351780 584960 351870
rect 428641 351386 428707 351389
rect 425194 351384 428707 351386
rect 425194 351328 428646 351384
rect 428702 351328 428707 351384
rect 425194 351326 428707 351328
rect 425194 350829 425254 351326
rect 428641 351323 428707 351326
rect -960 345402 480 345492
rect 3693 345402 3759 345405
rect -960 345400 3759 345402
rect -960 345344 3698 345400
rect 3754 345344 3759 345400
rect -960 345342 3759 345344
rect -960 345252 480 345342
rect 3693 345339 3759 345342
rect 37641 344994 37707 344997
rect 37641 344992 40110 344994
rect 37641 344936 37646 344992
rect 37702 344936 40110 344992
rect 37641 344934 40110 344936
rect 37641 344931 37707 344934
rect 428733 341730 428799 341733
rect 425194 341728 428799 341730
rect 425194 341672 428738 341728
rect 428794 341672 428799 341728
rect 425194 341670 428799 341672
rect 425194 341094 425254 341670
rect 428733 341667 428799 341670
rect 580625 338602 580691 338605
rect 583520 338602 584960 338692
rect 580625 338600 584960 338602
rect 580625 338544 580630 338600
rect 580686 338544 584960 338600
rect 580625 338542 584960 338544
rect 580625 338539 580691 338542
rect 583520 338452 584960 338542
rect 37825 336018 37891 336021
rect 37825 336016 40110 336018
rect 37825 335960 37830 336016
rect 37886 335960 40110 336016
rect 37825 335958 40110 335960
rect 37825 335955 37891 335958
rect 40050 335392 40110 335958
rect -960 332346 480 332436
rect 2773 332346 2839 332349
rect -960 332344 2839 332346
rect -960 332288 2778 332344
rect 2834 332288 2839 332344
rect -960 332286 2839 332288
rect -960 332196 480 332286
rect 2773 332283 2839 332286
rect 428549 332074 428615 332077
rect 425194 332072 428615 332074
rect 425194 332016 428554 332072
rect 428610 332016 428615 332072
rect 425194 332014 428615 332016
rect 425194 331398 425254 332014
rect 428549 332011 428615 332014
rect 37549 326498 37615 326501
rect 37549 326496 40110 326498
rect 37549 326440 37554 326496
rect 37610 326440 40110 326496
rect 37549 326438 40110 326440
rect 37549 326435 37615 326438
rect 40050 325869 40110 326438
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect 428825 322282 428891 322285
rect 425194 322280 428891 322282
rect 425194 322224 428830 322280
rect 428886 322224 428891 322280
rect 425194 322222 428891 322224
rect 425194 321645 425254 322222
rect 428825 322219 428891 322222
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 37917 316978 37983 316981
rect 37917 316976 40110 316978
rect 37917 316920 37922 316976
rect 37978 316920 40110 316976
rect 37917 316918 40110 316920
rect 37917 316915 37983 316918
rect 40050 316346 40110 316918
rect 428733 312626 428799 312629
rect 425194 312624 428799 312626
rect 425194 312568 428738 312624
rect 428794 312568 428799 312624
rect 425194 312566 428799 312568
rect 425194 311968 425254 312566
rect 428733 312563 428799 312566
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 37365 307322 37431 307325
rect 37365 307320 40110 307322
rect 37365 307264 37370 307320
rect 37426 307264 40110 307320
rect 37365 307262 40110 307264
rect 37365 307259 37431 307262
rect 40050 306803 40110 307262
rect -960 306234 480 306324
rect 3601 306234 3667 306237
rect -960 306232 3667 306234
rect -960 306176 3606 306232
rect 3662 306176 3667 306232
rect -960 306174 3667 306176
rect -960 306084 480 306174
rect 3601 306171 3667 306174
rect 428457 302834 428523 302837
rect 425194 302832 428523 302834
rect 425194 302776 428462 302832
rect 428518 302776 428523 302832
rect 425194 302774 428523 302776
rect 425194 302234 425254 302774
rect 428457 302771 428523 302774
rect 580257 298754 580323 298757
rect 583520 298754 584960 298844
rect 580257 298752 584960 298754
rect 580257 298696 580262 298752
rect 580318 298696 584960 298752
rect 580257 298694 584960 298696
rect 580257 298691 580323 298694
rect 583520 298604 584960 298694
rect 37549 297666 37615 297669
rect 37549 297664 40110 297666
rect 37549 297608 37554 297664
rect 37610 297608 40110 297664
rect 37549 297606 40110 297608
rect 37549 297603 37615 297606
rect 40050 297280 40110 297606
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 425194 292498 425254 292518
rect 428457 292498 428523 292501
rect 425194 292496 428523 292498
rect 425194 292440 428462 292496
rect 428518 292440 428523 292496
rect 425194 292438 428523 292440
rect 428457 292435 428523 292438
rect 37733 288282 37799 288285
rect 37733 288280 40110 288282
rect 37733 288224 37738 288280
rect 37794 288224 40110 288280
rect 37733 288222 40110 288224
rect 37733 288219 37799 288222
rect 40050 287776 40110 288222
rect 580349 285426 580415 285429
rect 583520 285426 584960 285516
rect 580349 285424 584960 285426
rect 580349 285368 580354 285424
rect 580410 285368 584960 285424
rect 580349 285366 584960 285368
rect 580349 285363 580415 285366
rect 583520 285276 584960 285366
rect 429009 282842 429075 282845
rect 425194 282840 429075 282842
rect 425194 282784 429014 282840
rect 429070 282784 429075 282840
rect 425194 282782 429075 282784
rect 429009 282779 429075 282782
rect -960 280122 480 280212
rect 3693 280122 3759 280125
rect -960 280120 3759 280122
rect -960 280064 3698 280120
rect 3754 280064 3759 280120
rect -960 280062 3759 280064
rect -960 279972 480 280062
rect 3693 280059 3759 280062
rect 37733 278490 37799 278493
rect 37733 278488 40110 278490
rect 37733 278432 37738 278488
rect 37794 278432 40110 278488
rect 37733 278430 40110 278432
rect 37733 278427 37799 278430
rect 40050 278234 40110 278430
rect 428549 273186 428615 273189
rect 425194 273184 428615 273186
rect 425194 273128 428554 273184
rect 428610 273128 428615 273184
rect 425194 273126 428615 273128
rect 425194 273107 425254 273126
rect 428549 273123 428615 273126
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect 37917 268970 37983 268973
rect 37917 268968 40110 268970
rect 37917 268912 37922 268968
rect 37978 268912 40110 268968
rect 37917 268910 40110 268912
rect 37917 268907 37983 268910
rect 40050 268730 40110 268910
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 428641 263530 428707 263533
rect 425194 263528 428707 263530
rect 425194 263472 428646 263528
rect 428702 263472 428707 263528
rect 425194 263470 428707 263472
rect 425194 263373 425254 263470
rect 428641 263467 428707 263470
rect 37365 258090 37431 258093
rect 37365 258088 37474 258090
rect 37365 258032 37370 258088
rect 37426 258032 37474 258088
rect 37365 258027 37474 258032
rect 37414 257954 37474 258027
rect 40050 257954 40110 259187
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect 37414 257894 40110 257954
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 428917 253874 428983 253877
rect 425194 253872 428983 253874
rect 425194 253816 428922 253872
rect 428978 253816 428983 253872
rect 425194 253814 428983 253816
rect 425194 253658 425254 253814
rect 428917 253811 428983 253814
rect 37917 249658 37983 249661
rect 37917 249656 39498 249658
rect 37917 249600 37922 249656
rect 37978 249600 40020 249656
rect 37917 249598 40020 249600
rect 37917 249595 37983 249598
rect 39438 249596 40020 249598
rect 579797 245578 579863 245581
rect 583520 245578 584960 245668
rect 579797 245576 584960 245578
rect 579797 245520 579802 245576
rect 579858 245520 584960 245576
rect 579797 245518 584960 245520
rect 579797 245515 579863 245518
rect 583520 245428 584960 245518
rect 428641 244218 428707 244221
rect 425194 244216 428707 244218
rect 425194 244160 428646 244216
rect 428702 244160 428707 244216
rect 425194 244158 428707 244160
rect 425194 243962 425254 244158
rect 428641 244155 428707 244158
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 37365 240138 37431 240141
rect 37365 240136 39498 240138
rect 37365 240080 37370 240136
rect 37426 240113 39498 240136
rect 37426 240080 40020 240113
rect 37365 240078 40020 240080
rect 37365 240075 37431 240078
rect 39438 240053 40020 240078
rect 428457 234562 428523 234565
rect 425194 234560 428523 234562
rect 425194 234504 428462 234560
rect 428518 234504 428523 234560
rect 425194 234502 428523 234504
rect 425194 234227 425254 234502
rect 428457 234499 428523 234502
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 37641 230618 37707 230621
rect 37641 230616 39498 230618
rect 37641 230560 37646 230616
rect 37702 230590 39498 230616
rect 37702 230560 40020 230590
rect 37641 230558 40020 230560
rect 37641 230555 37707 230558
rect 39438 230530 40020 230558
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 428549 224906 428615 224909
rect 425194 224904 428615 224906
rect 425194 224848 428554 224904
rect 428610 224848 428615 224904
rect 425194 224846 428615 224848
rect 425194 224512 425254 224846
rect 428549 224843 428615 224846
rect 37733 221642 37799 221645
rect 37733 221640 40110 221642
rect 37733 221584 37738 221640
rect 37794 221584 40110 221640
rect 37733 221582 40110 221584
rect 37733 221579 37799 221582
rect 40050 221018 40110 221582
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 428641 215250 428707 215253
rect 425194 215248 428707 215250
rect 425194 215192 428646 215248
rect 428702 215192 428707 215248
rect 425194 215190 428707 215192
rect -960 214978 480 215068
rect 3601 214978 3667 214981
rect -960 214976 3667 214978
rect -960 214920 3606 214976
rect 3662 214920 3667 214976
rect -960 214918 3667 214920
rect -960 214828 480 214918
rect 3601 214915 3667 214918
rect 425194 214816 425254 215190
rect 428641 215187 428707 215190
rect 37825 212122 37891 212125
rect 37825 212120 40110 212122
rect 37825 212064 37830 212120
rect 37886 212064 40110 212120
rect 37825 212062 40110 212064
rect 37825 212059 37891 212062
rect 40050 211494 40110 212062
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 428457 205594 428523 205597
rect 425194 205592 428523 205594
rect 425194 205536 428462 205592
rect 428518 205536 428523 205592
rect 583520 205580 584960 205670
rect 425194 205534 428523 205536
rect 425194 205101 425254 205534
rect 428457 205531 428523 205534
rect 37733 202602 37799 202605
rect 37733 202600 40110 202602
rect 37733 202544 37738 202600
rect 37794 202544 40110 202600
rect 37733 202542 40110 202544
rect 37733 202539 37799 202542
rect -960 201922 480 202012
rect 40050 201952 40110 202542
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 428549 195938 428615 195941
rect 425194 195936 428615 195938
rect 425194 195880 428554 195936
rect 428610 195880 428615 195936
rect 425194 195878 428615 195880
rect 425194 195366 425254 195878
rect 428549 195875 428615 195878
rect 37733 192946 37799 192949
rect 37733 192944 40110 192946
rect 37733 192888 37738 192944
rect 37794 192888 40110 192944
rect 37733 192886 40110 192888
rect 37733 192883 37799 192886
rect 40050 192429 40110 192886
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 428641 186282 428707 186285
rect 425194 186280 428707 186282
rect 425194 186224 428646 186280
rect 428702 186224 428707 186280
rect 425194 186222 428707 186224
rect 425194 185690 425254 186222
rect 428641 186219 428707 186222
rect 37917 183426 37983 183429
rect 37917 183424 40110 183426
rect 37917 183368 37922 183424
rect 37978 183368 40110 183424
rect 37917 183366 40110 183368
rect 37917 183363 37983 183366
rect 40050 182925 40110 183366
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 428457 176626 428523 176629
rect 425194 176624 428523 176626
rect 425194 176568 428462 176624
rect 428518 176568 428523 176624
rect 425194 176566 428523 176568
rect -960 175946 480 176036
rect 425194 175955 425254 176566
rect 428457 176563 428523 176566
rect 3509 175946 3575 175949
rect -960 175944 3575 175946
rect -960 175888 3514 175944
rect 3570 175888 3575 175944
rect -960 175886 3575 175888
rect -960 175796 480 175886
rect 3509 175883 3575 175886
rect 37733 173634 37799 173637
rect 37733 173632 40110 173634
rect 37733 173576 37738 173632
rect 37794 173576 40110 173632
rect 37733 173574 40110 173576
rect 37733 173571 37799 173574
rect 40050 173402 40110 173574
rect 428549 166834 428615 166837
rect 425194 166832 428615 166834
rect 425194 166776 428554 166832
rect 428610 166776 428615 166832
rect 425194 166774 428615 166776
rect 425194 166240 425254 166774
rect 428549 166771 428615 166774
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 37917 164114 37983 164117
rect 37917 164112 40110 164114
rect 37917 164056 37922 164112
rect 37978 164056 40110 164112
rect 37917 164054 40110 164056
rect 37917 164051 37983 164054
rect 40050 163859 40110 164054
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 428457 157178 428523 157181
rect 425194 157176 428523 157178
rect 425194 157120 428462 157176
rect 428518 157120 428523 157176
rect 425194 157118 428523 157120
rect 425194 156525 425254 157118
rect 428457 157115 428523 157118
rect 37641 154322 37707 154325
rect 40050 154322 40110 154336
rect 37641 154320 40110 154322
rect 37641 154264 37646 154320
rect 37702 154264 40110 154320
rect 37641 154262 40110 154264
rect 37641 154259 37707 154262
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 429101 147386 429167 147389
rect 425194 147384 429167 147386
rect 425194 147328 429106 147384
rect 429162 147328 429167 147384
rect 425194 147326 429167 147328
rect 425194 146810 425254 147326
rect 429101 147323 429167 147326
rect 37917 144802 37983 144805
rect 39438 144802 40020 144824
rect 37917 144800 40020 144802
rect 37917 144744 37922 144800
rect 37978 144764 40020 144800
rect 37978 144744 39498 144764
rect 37917 144742 39498 144744
rect 37917 144739 37983 144742
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 428825 137594 428891 137597
rect 425194 137592 428891 137594
rect 425194 137536 428830 137592
rect 428886 137536 428891 137592
rect 425194 137534 428891 137536
rect 425194 137075 425254 137534
rect 428825 137531 428891 137534
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 37549 135826 37615 135829
rect 37549 135824 40110 135826
rect 37549 135768 37554 135824
rect 37610 135768 40110 135824
rect 37549 135766 40110 135768
rect 37549 135763 37615 135766
rect 40050 135232 40110 135766
rect 425194 127122 425254 127379
rect 428917 127122 428983 127125
rect 425194 127120 428983 127122
rect 425194 127064 428922 127120
rect 428978 127064 428983 127120
rect 425194 127062 428983 127064
rect 428917 127059 428983 127062
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 37733 125762 37799 125765
rect 37733 125760 39498 125762
rect 37733 125704 37738 125760
rect 37794 125758 39498 125760
rect 37794 125704 40020 125758
rect 37733 125702 40020 125704
rect 37733 125699 37799 125702
rect 39438 125698 40020 125702
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 425194 117330 425254 117645
rect 428457 117330 428523 117333
rect 425194 117328 428523 117330
rect 425194 117272 428462 117328
rect 428518 117272 428523 117328
rect 425194 117270 428523 117272
rect 428457 117267 428523 117270
rect 37917 115970 37983 115973
rect 40050 115970 40110 116186
rect 37917 115968 40110 115970
rect 37917 115912 37922 115968
rect 37978 115912 40110 115968
rect 37917 115910 40110 115912
rect 37917 115907 37983 115910
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 425194 107674 425254 107930
rect 428457 107674 428523 107677
rect 425194 107672 428523 107674
rect 425194 107616 428462 107672
rect 428518 107616 428523 107672
rect 425194 107614 428523 107616
rect 428457 107611 428523 107614
rect 37917 106314 37983 106317
rect 40050 106314 40110 106662
rect 37917 106312 40110 106314
rect 37917 106256 37922 106312
rect 37978 106256 40110 106312
rect 37917 106254 40110 106256
rect 37917 106251 37983 106254
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 425194 98018 425254 98253
rect 428549 98018 428615 98021
rect 425194 98016 428615 98018
rect 425194 97960 428554 98016
rect 428610 97960 428615 98016
rect 425194 97958 428615 97960
rect 428549 97955 428615 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 38009 96658 38075 96661
rect 40050 96658 40110 97120
rect 38009 96656 40110 96658
rect 38009 96600 38014 96656
rect 38070 96600 40110 96656
rect 38009 96598 40110 96600
rect 38009 96595 38075 96598
rect 425194 88362 425254 88499
rect 428457 88362 428523 88365
rect 425194 88360 428523 88362
rect 425194 88304 428462 88360
rect 428518 88304 428523 88360
rect 425194 88302 428523 88304
rect 428457 88299 428523 88302
rect 37917 87002 37983 87005
rect 40050 87002 40110 87597
rect 37917 87000 40110 87002
rect 37917 86944 37922 87000
rect 37978 86944 40110 87000
rect 37917 86942 40110 86944
rect 37917 86939 37983 86942
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 425194 78706 425254 78803
rect 428549 78706 428615 78709
rect 425194 78704 428615 78706
rect 425194 78648 428554 78704
rect 428610 78648 428615 78704
rect 425194 78646 428615 78648
rect 428549 78643 428615 78646
rect 38009 77482 38075 77485
rect 40050 77482 40110 78054
rect 38009 77480 40110 77482
rect 38009 77424 38014 77480
rect 38070 77424 40110 77480
rect 38009 77422 40110 77424
rect 38009 77419 38075 77422
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 428457 69186 428523 69189
rect 425194 69184 428523 69186
rect 425194 69128 428462 69184
rect 428518 69128 428523 69184
rect 425194 69126 428523 69128
rect 425194 69107 425254 69126
rect 428457 69123 428523 69126
rect 37917 67962 37983 67965
rect 40050 67962 40110 68531
rect 37917 67960 40110 67962
rect 37917 67904 37922 67960
rect 37978 67904 40110 67960
rect 37917 67902 40110 67904
rect 37917 67899 37983 67902
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect 428641 59394 428707 59397
rect 425194 59392 428707 59394
rect 425194 59336 428646 59392
rect 428702 59336 428707 59392
rect 425194 59334 428707 59336
rect 428641 59331 428707 59334
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 38101 58442 38167 58445
rect 40050 58442 40110 59008
rect 38101 58440 40110 58442
rect 38101 58384 38106 58440
rect 38162 58384 40110 58440
rect 38101 58382 40110 58384
rect 38101 58379 38167 58382
rect 38009 49330 38075 49333
rect 38009 49328 39498 49330
rect 38009 49272 38014 49328
rect 38070 49322 39498 49328
rect 38070 49272 40020 49322
rect 38009 49270 40020 49272
rect 38009 49267 38075 49270
rect 39438 49262 40020 49270
rect 425194 49058 425254 49619
rect 428549 49058 428615 49061
rect 425194 49056 428615 49058
rect 425194 49000 428554 49056
rect 428610 49000 428615 49056
rect 425194 48998 428615 49000
rect 428549 48995 428615 48998
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 37917 40218 37983 40221
rect 37917 40216 40110 40218
rect 37917 40160 37922 40216
rect 37978 40160 40110 40216
rect 37917 40158 40110 40160
rect 37917 40155 37983 40158
rect 40050 40154 40110 40158
rect 425194 40082 425254 40403
rect 428457 40082 428523 40085
rect 425194 40080 428523 40082
rect 425194 40024 428462 40080
rect 428518 40024 428523 40080
rect 425194 40022 428523 40024
rect 428457 40019 428523 40022
rect 579889 33146 579955 33149
rect 583520 33146 584960 33236
rect 579889 33144 584960 33146
rect 579889 33088 579894 33144
rect 579950 33088 584960 33144
rect 579889 33086 584960 33088
rect 579889 33083 579955 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 579889 19818 579955 19821
rect 583520 19818 584960 19908
rect 579889 19816 584960 19818
rect 579889 19760 579894 19816
rect 579950 19760 584960 19816
rect 579889 19758 584960 19760
rect 579889 19755 579955 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 5257 3362 5323 3365
rect 120257 3362 120323 3365
rect 5257 3360 120323 3362
rect 5257 3304 5262 3360
rect 5318 3304 120262 3360
rect 120318 3304 120323 3360
rect 5257 3302 120323 3304
rect 5257 3299 5323 3302
rect 120257 3299 120323 3302
rect 305545 3362 305611 3365
rect 361573 3362 361639 3365
rect 305545 3360 361639 3362
rect 305545 3304 305550 3360
rect 305606 3304 361578 3360
rect 361634 3304 361639 3360
rect 305545 3302 361639 3304
rect 305545 3299 305611 3302
rect 361573 3299 361639 3302
rect 398833 3362 398899 3365
rect 479333 3362 479399 3365
rect 398833 3360 479399 3362
rect 398833 3304 398838 3360
rect 398894 3304 479338 3360
rect 479394 3304 479399 3360
rect 398833 3302 479399 3304
rect 398833 3299 398899 3302
rect 479333 3299 479399 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 561044 38414 578898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 561044 42134 582618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 561044 45854 586338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 561044 49574 590058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561044 56414 596898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 561044 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 561044 63854 568338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 561044 67574 572058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 561044 74414 578898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 561044 78134 582618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 561044 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 561044 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561044 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 561044 96134 564618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 561044 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 561044 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 561044 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 561044 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 561044 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 561044 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561044 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 561044 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 561044 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 561044 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 561044 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 561044 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 561044 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 561044 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561044 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 561044 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 561044 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 561044 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 561044 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 561044 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 561044 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 561044 193574 590058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561044 200414 596898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 561044 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 561044 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 561044 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 561044 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 561044 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 561044 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 561044 229574 590058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561044 236414 596898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 561044 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 561044 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 561044 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 561044 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 561044 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 561044 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 561044 265574 590058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561044 272414 596898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 561044 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 561044 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 561044 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 561044 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 561044 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 561044 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 561044 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561044 308414 596898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 561044 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 561044 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 561044 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 561044 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 561044 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 561044 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 561044 337574 590058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561044 344414 596898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 561044 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 561044 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 561044 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 561044 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 561044 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 561044 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 561044 373574 590058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561044 380414 596898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 561044 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 561044 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 561044 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 561044 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 561044 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 561044 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 561044 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561044 416414 596898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 561044 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 561044 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 561044 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 42556 543454 43356 543486
rect 42556 543218 42678 543454
rect 42914 543218 42998 543454
rect 43234 543218 43356 543454
rect 42556 543134 43356 543218
rect 42556 542898 42678 543134
rect 42914 542898 42998 543134
rect 43234 542898 43356 543134
rect 42556 542866 43356 542898
rect 200527 543454 200927 543486
rect 200527 543218 200609 543454
rect 200845 543218 200927 543454
rect 200527 543134 200927 543218
rect 200527 542898 200609 543134
rect 200845 542898 200927 543134
rect 200527 542866 200927 542898
rect 416915 543454 417315 543486
rect 416915 543218 416997 543454
rect 417233 543218 417315 543454
rect 416915 543134 417315 543218
rect 416915 542898 416997 543134
rect 417233 542898 417315 543134
rect 416915 542866 417315 542898
rect 421940 543454 422740 543486
rect 421940 543218 422062 543454
rect 422298 543218 422382 543454
rect 422618 543218 422740 543454
rect 421940 543134 422740 543218
rect 421940 542898 422062 543134
rect 422298 542898 422382 543134
rect 422618 542898 422740 543134
rect 421940 542866 422740 542898
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 41396 525454 42196 525486
rect 41396 525218 41518 525454
rect 41754 525218 41838 525454
rect 42074 525218 42196 525454
rect 41396 525134 42196 525218
rect 41396 524898 41518 525134
rect 41754 524898 41838 525134
rect 42074 524898 42196 525134
rect 41396 524866 42196 524898
rect 199767 525454 200167 525486
rect 199767 525218 199849 525454
rect 200085 525218 200167 525454
rect 199767 525134 200167 525218
rect 199767 524898 199849 525134
rect 200085 524898 200167 525134
rect 199767 524866 200167 524898
rect 204981 525454 205329 525486
rect 204981 525218 205037 525454
rect 205273 525218 205329 525454
rect 204981 525134 205329 525218
rect 204981 524898 205037 525134
rect 205273 524898 205329 525134
rect 204981 524866 205329 524898
rect 300045 525454 300393 525486
rect 300045 525218 300101 525454
rect 300337 525218 300393 525454
rect 300045 525134 300393 525218
rect 300045 524898 300101 525134
rect 300337 524898 300393 525134
rect 300045 524866 300393 524898
rect 317409 525454 317757 525486
rect 317409 525218 317465 525454
rect 317701 525218 317757 525454
rect 317409 525134 317757 525218
rect 317409 524898 317465 525134
rect 317701 524898 317757 525134
rect 317409 524866 317757 524898
rect 412473 525454 412821 525486
rect 412473 525218 412529 525454
rect 412765 525218 412821 525454
rect 412473 525134 412821 525218
rect 412473 524898 412529 525134
rect 412765 524898 412821 525134
rect 412473 524866 412821 524898
rect 417675 525454 418075 525486
rect 417675 525218 417757 525454
rect 417993 525218 418075 525454
rect 417675 525134 418075 525218
rect 417675 524898 417757 525134
rect 417993 524898 418075 525134
rect 417675 524866 418075 524898
rect 423100 525454 423900 525486
rect 423100 525218 423222 525454
rect 423458 525218 423542 525454
rect 423778 525218 423900 525454
rect 423100 525134 423900 525218
rect 423100 524898 423222 525134
rect 423458 524898 423542 525134
rect 423778 524898 423900 525134
rect 423100 524866 423900 524898
rect 42556 507454 43356 507486
rect 42556 507218 42678 507454
rect 42914 507218 42998 507454
rect 43234 507218 43356 507454
rect 42556 507134 43356 507218
rect 42556 506898 42678 507134
rect 42914 506898 42998 507134
rect 43234 506898 43356 507134
rect 42556 506866 43356 506898
rect 200527 507454 200927 507486
rect 200527 507218 200609 507454
rect 200845 507218 200927 507454
rect 200527 507134 200927 507218
rect 200527 506898 200609 507134
rect 200845 506898 200927 507134
rect 200527 506866 200927 506898
rect 205661 507454 206009 507486
rect 205661 507218 205717 507454
rect 205953 507218 206009 507454
rect 205661 507134 206009 507218
rect 205661 506898 205717 507134
rect 205953 506898 206009 507134
rect 205661 506866 206009 506898
rect 299365 507454 299713 507486
rect 299365 507218 299421 507454
rect 299657 507218 299713 507454
rect 299365 507134 299713 507218
rect 299365 506898 299421 507134
rect 299657 506898 299713 507134
rect 299365 506866 299713 506898
rect 318089 507454 318437 507486
rect 318089 507218 318145 507454
rect 318381 507218 318437 507454
rect 318089 507134 318437 507218
rect 318089 506898 318145 507134
rect 318381 506898 318437 507134
rect 318089 506866 318437 506898
rect 411793 507454 412141 507486
rect 411793 507218 411849 507454
rect 412085 507218 412141 507454
rect 411793 507134 412141 507218
rect 411793 506898 411849 507134
rect 412085 506898 412141 507134
rect 411793 506866 412141 506898
rect 416915 507454 417315 507486
rect 416915 507218 416997 507454
rect 417233 507218 417315 507454
rect 416915 507134 417315 507218
rect 416915 506898 416997 507134
rect 417233 506898 417315 507134
rect 416915 506866 417315 506898
rect 421940 507454 422740 507486
rect 421940 507218 422062 507454
rect 422298 507218 422382 507454
rect 422618 507218 422740 507454
rect 421940 507134 422740 507218
rect 421940 506898 422062 507134
rect 422298 506898 422382 507134
rect 422618 506898 422740 507134
rect 421940 506866 422740 506898
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 41396 489454 42196 489486
rect 41396 489218 41518 489454
rect 41754 489218 41838 489454
rect 42074 489218 42196 489454
rect 41396 489134 42196 489218
rect 41396 488898 41518 489134
rect 41754 488898 41838 489134
rect 42074 488898 42196 489134
rect 41396 488866 42196 488898
rect 199767 489454 200167 489486
rect 199767 489218 199849 489454
rect 200085 489218 200167 489454
rect 199767 489134 200167 489218
rect 199767 488898 199849 489134
rect 200085 488898 200167 489134
rect 199767 488866 200167 488898
rect 204981 489454 205329 489486
rect 204981 489218 205037 489454
rect 205273 489218 205329 489454
rect 204981 489134 205329 489218
rect 204981 488898 205037 489134
rect 205273 488898 205329 489134
rect 204981 488866 205329 488898
rect 300045 489454 300393 489486
rect 300045 489218 300101 489454
rect 300337 489218 300393 489454
rect 300045 489134 300393 489218
rect 300045 488898 300101 489134
rect 300337 488898 300393 489134
rect 300045 488866 300393 488898
rect 317409 489454 317757 489486
rect 317409 489218 317465 489454
rect 317701 489218 317757 489454
rect 317409 489134 317757 489218
rect 317409 488898 317465 489134
rect 317701 488898 317757 489134
rect 317409 488866 317757 488898
rect 412473 489454 412821 489486
rect 412473 489218 412529 489454
rect 412765 489218 412821 489454
rect 412473 489134 412821 489218
rect 412473 488898 412529 489134
rect 412765 488898 412821 489134
rect 412473 488866 412821 488898
rect 417675 489454 418075 489486
rect 417675 489218 417757 489454
rect 417993 489218 418075 489454
rect 417675 489134 418075 489218
rect 417675 488898 417757 489134
rect 417993 488898 418075 489134
rect 417675 488866 418075 488898
rect 423100 489454 423900 489486
rect 423100 489218 423222 489454
rect 423458 489218 423542 489454
rect 423778 489218 423900 489454
rect 423100 489134 423900 489218
rect 423100 488898 423222 489134
rect 423458 488898 423542 489134
rect 423778 488898 423900 489134
rect 423100 488866 423900 488898
rect 42556 471454 43356 471486
rect 42556 471218 42678 471454
rect 42914 471218 42998 471454
rect 43234 471218 43356 471454
rect 42556 471134 43356 471218
rect 42556 470898 42678 471134
rect 42914 470898 42998 471134
rect 43234 470898 43356 471134
rect 42556 470866 43356 470898
rect 200527 471454 200927 471486
rect 200527 471218 200609 471454
rect 200845 471218 200927 471454
rect 200527 471134 200927 471218
rect 200527 470898 200609 471134
rect 200845 470898 200927 471134
rect 200527 470866 200927 470898
rect 205661 471454 206009 471486
rect 205661 471218 205717 471454
rect 205953 471218 206009 471454
rect 205661 471134 206009 471218
rect 205661 470898 205717 471134
rect 205953 470898 206009 471134
rect 205661 470866 206009 470898
rect 299365 471454 299713 471486
rect 299365 471218 299421 471454
rect 299657 471218 299713 471454
rect 299365 471134 299713 471218
rect 299365 470898 299421 471134
rect 299657 470898 299713 471134
rect 299365 470866 299713 470898
rect 318089 471454 318437 471486
rect 318089 471218 318145 471454
rect 318381 471218 318437 471454
rect 318089 471134 318437 471218
rect 318089 470898 318145 471134
rect 318381 470898 318437 471134
rect 318089 470866 318437 470898
rect 411793 471454 412141 471486
rect 411793 471218 411849 471454
rect 412085 471218 412141 471454
rect 411793 471134 412141 471218
rect 411793 470898 411849 471134
rect 412085 470898 412141 471134
rect 411793 470866 412141 470898
rect 416915 471454 417315 471486
rect 416915 471218 416997 471454
rect 417233 471218 417315 471454
rect 416915 471134 417315 471218
rect 416915 470898 416997 471134
rect 417233 470898 417315 471134
rect 416915 470866 417315 470898
rect 421940 471454 422740 471486
rect 421940 471218 422062 471454
rect 422298 471218 422382 471454
rect 422618 471218 422740 471454
rect 421940 471134 422740 471218
rect 421940 470898 422062 471134
rect 422298 470898 422382 471134
rect 422618 470898 422740 471134
rect 421940 470866 422740 470898
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 41396 453454 42196 453486
rect 41396 453218 41518 453454
rect 41754 453218 41838 453454
rect 42074 453218 42196 453454
rect 41396 453134 42196 453218
rect 41396 452898 41518 453134
rect 41754 452898 41838 453134
rect 42074 452898 42196 453134
rect 41396 452866 42196 452898
rect 423100 453454 423900 453486
rect 423100 453218 423222 453454
rect 423458 453218 423542 453454
rect 423778 453218 423900 453454
rect 423100 453134 423900 453218
rect 423100 452898 423222 453134
rect 423458 452898 423542 453134
rect 423778 452898 423900 453134
rect 423100 452866 423900 452898
rect 42556 435454 43356 435486
rect 42556 435218 42678 435454
rect 42914 435218 42998 435454
rect 43234 435218 43356 435454
rect 42556 435134 43356 435218
rect 42556 434898 42678 435134
rect 42914 434898 42998 435134
rect 43234 434898 43356 435134
rect 42556 434866 43356 434898
rect 198552 435454 198900 435486
rect 198552 435218 198608 435454
rect 198844 435218 198900 435454
rect 198552 435134 198900 435218
rect 198552 434898 198608 435134
rect 198844 434898 198900 435134
rect 198552 434866 198900 434898
rect 292256 435454 292604 435486
rect 292256 435218 292312 435454
rect 292548 435218 292604 435454
rect 292256 435134 292604 435218
rect 292256 434898 292312 435134
rect 292548 434898 292604 435134
rect 292256 434866 292604 434898
rect 325108 435454 325456 435486
rect 325108 435218 325164 435454
rect 325400 435218 325456 435454
rect 325108 435134 325456 435218
rect 325108 434898 325164 435134
rect 325400 434898 325456 435134
rect 325108 434866 325456 434898
rect 418812 435454 419160 435486
rect 418812 435218 418868 435454
rect 419104 435218 419160 435454
rect 418812 435134 419160 435218
rect 418812 434898 418868 435134
rect 419104 434898 419160 435134
rect 418812 434866 419160 434898
rect 421940 435454 422740 435486
rect 421940 435218 422062 435454
rect 422298 435218 422382 435454
rect 422618 435218 422740 435454
rect 421940 435134 422740 435218
rect 421940 434898 422062 435134
rect 422298 434898 422382 435134
rect 422618 434898 422740 435134
rect 421940 434866 422740 434898
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 41396 417454 42196 417486
rect 41396 417218 41518 417454
rect 41754 417218 41838 417454
rect 42074 417218 42196 417454
rect 41396 417134 42196 417218
rect 41396 416898 41518 417134
rect 41754 416898 41838 417134
rect 42074 416898 42196 417134
rect 41396 416866 42196 416898
rect 197872 417454 198220 417486
rect 197872 417218 197928 417454
rect 198164 417218 198220 417454
rect 197872 417134 198220 417218
rect 197872 416898 197928 417134
rect 198164 416898 198220 417134
rect 197872 416866 198220 416898
rect 292936 417454 293284 417486
rect 292936 417218 292992 417454
rect 293228 417218 293284 417454
rect 292936 417134 293284 417218
rect 292936 416898 292992 417134
rect 293228 416898 293284 417134
rect 292936 416866 293284 416898
rect 324428 417454 324776 417486
rect 324428 417218 324484 417454
rect 324720 417218 324776 417454
rect 324428 417134 324776 417218
rect 324428 416898 324484 417134
rect 324720 416898 324776 417134
rect 324428 416866 324776 416898
rect 419492 417454 419840 417486
rect 419492 417218 419548 417454
rect 419784 417218 419840 417454
rect 419492 417134 419840 417218
rect 419492 416898 419548 417134
rect 419784 416898 419840 417134
rect 419492 416866 419840 416898
rect 423100 417454 423900 417486
rect 423100 417218 423222 417454
rect 423458 417218 423542 417454
rect 423778 417218 423900 417454
rect 423100 417134 423900 417218
rect 423100 416898 423222 417134
rect 423458 416898 423542 417134
rect 423778 416898 423900 417134
rect 423100 416866 423900 416898
rect 42556 399454 43356 399486
rect 42556 399218 42678 399454
rect 42914 399218 42998 399454
rect 43234 399218 43356 399454
rect 42556 399134 43356 399218
rect 42556 398898 42678 399134
rect 42914 398898 42998 399134
rect 43234 398898 43356 399134
rect 42556 398866 43356 398898
rect 198552 399454 198900 399486
rect 198552 399218 198608 399454
rect 198844 399218 198900 399454
rect 198552 399134 198900 399218
rect 198552 398898 198608 399134
rect 198844 398898 198900 399134
rect 198552 398866 198900 398898
rect 292256 399454 292604 399486
rect 292256 399218 292312 399454
rect 292548 399218 292604 399454
rect 292256 399134 292604 399218
rect 292256 398898 292312 399134
rect 292548 398898 292604 399134
rect 292256 398866 292604 398898
rect 325108 399454 325456 399486
rect 325108 399218 325164 399454
rect 325400 399218 325456 399454
rect 325108 399134 325456 399218
rect 325108 398898 325164 399134
rect 325400 398898 325456 399134
rect 325108 398866 325456 398898
rect 418812 399454 419160 399486
rect 418812 399218 418868 399454
rect 419104 399218 419160 399454
rect 418812 399134 419160 399218
rect 418812 398898 418868 399134
rect 419104 398898 419160 399134
rect 418812 398866 419160 398898
rect 421940 399454 422740 399486
rect 421940 399218 422062 399454
rect 422298 399218 422382 399454
rect 422618 399218 422740 399454
rect 421940 399134 422740 399218
rect 421940 398898 422062 399134
rect 422298 398898 422382 399134
rect 422618 398898 422740 399134
rect 421940 398866 422740 398898
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 41396 381454 42196 381486
rect 41396 381218 41518 381454
rect 41754 381218 41838 381454
rect 42074 381218 42196 381454
rect 41396 381134 42196 381218
rect 41396 380898 41518 381134
rect 41754 380898 41838 381134
rect 42074 380898 42196 381134
rect 41396 380866 42196 380898
rect 197872 381454 198220 381486
rect 197872 381218 197928 381454
rect 198164 381218 198220 381454
rect 197872 381134 198220 381218
rect 197872 380898 197928 381134
rect 198164 380898 198220 381134
rect 197872 380866 198220 380898
rect 292936 381454 293284 381486
rect 292936 381218 292992 381454
rect 293228 381218 293284 381454
rect 292936 381134 293284 381218
rect 292936 380898 292992 381134
rect 293228 380898 293284 381134
rect 292936 380866 293284 380898
rect 324428 381454 324776 381486
rect 324428 381218 324484 381454
rect 324720 381218 324776 381454
rect 324428 381134 324776 381218
rect 324428 380898 324484 381134
rect 324720 380898 324776 381134
rect 324428 380866 324776 380898
rect 419492 381454 419840 381486
rect 419492 381218 419548 381454
rect 419784 381218 419840 381454
rect 419492 381134 419840 381218
rect 419492 380898 419548 381134
rect 419784 380898 419840 381134
rect 419492 380866 419840 380898
rect 423100 381454 423900 381486
rect 423100 381218 423222 381454
rect 423458 381218 423542 381454
rect 423778 381218 423900 381454
rect 423100 381134 423900 381218
rect 423100 380898 423222 381134
rect 423458 380898 423542 381134
rect 423778 380898 423900 381134
rect 423100 380866 423900 380898
rect 42556 363454 43356 363486
rect 42556 363218 42678 363454
rect 42914 363218 42998 363454
rect 43234 363218 43356 363454
rect 42556 363134 43356 363218
rect 42556 362898 42678 363134
rect 42914 362898 42998 363134
rect 43234 362898 43356 363134
rect 42556 362866 43356 362898
rect 421940 363454 422740 363486
rect 421940 363218 422062 363454
rect 422298 363218 422382 363454
rect 422618 363218 422740 363454
rect 421940 363134 422740 363218
rect 421940 362898 422062 363134
rect 422298 362898 422382 363134
rect 422618 362898 422740 363134
rect 421940 362866 422740 362898
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 41396 345454 42196 345486
rect 41396 345218 41518 345454
rect 41754 345218 41838 345454
rect 42074 345218 42196 345454
rect 41396 345134 42196 345218
rect 41396 344898 41518 345134
rect 41754 344898 41838 345134
rect 42074 344898 42196 345134
rect 41396 344866 42196 344898
rect 423100 345454 423900 345486
rect 423100 345218 423222 345454
rect 423458 345218 423542 345454
rect 423778 345218 423900 345454
rect 423100 345134 423900 345218
rect 423100 344898 423222 345134
rect 423458 344898 423542 345134
rect 423778 344898 423900 345134
rect 423100 344866 423900 344898
rect 42556 327454 43356 327486
rect 42556 327218 42678 327454
rect 42914 327218 42998 327454
rect 43234 327218 43356 327454
rect 42556 327134 43356 327218
rect 42556 326898 42678 327134
rect 42914 326898 42998 327134
rect 43234 326898 43356 327134
rect 42556 326866 43356 326898
rect 198552 327454 198900 327486
rect 198552 327218 198608 327454
rect 198844 327218 198900 327454
rect 198552 327134 198900 327218
rect 198552 326898 198608 327134
rect 198844 326898 198900 327134
rect 198552 326866 198900 326898
rect 292256 327454 292604 327486
rect 292256 327218 292312 327454
rect 292548 327218 292604 327454
rect 292256 327134 292604 327218
rect 292256 326898 292312 327134
rect 292548 326898 292604 327134
rect 292256 326866 292604 326898
rect 325108 327454 325456 327486
rect 325108 327218 325164 327454
rect 325400 327218 325456 327454
rect 325108 327134 325456 327218
rect 325108 326898 325164 327134
rect 325400 326898 325456 327134
rect 325108 326866 325456 326898
rect 418812 327454 419160 327486
rect 418812 327218 418868 327454
rect 419104 327218 419160 327454
rect 418812 327134 419160 327218
rect 418812 326898 418868 327134
rect 419104 326898 419160 327134
rect 418812 326866 419160 326898
rect 421940 327454 422740 327486
rect 421940 327218 422062 327454
rect 422298 327218 422382 327454
rect 422618 327218 422740 327454
rect 421940 327134 422740 327218
rect 421940 326898 422062 327134
rect 422298 326898 422382 327134
rect 422618 326898 422740 327134
rect 421940 326866 422740 326898
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 41396 309454 42196 309486
rect 41396 309218 41518 309454
rect 41754 309218 41838 309454
rect 42074 309218 42196 309454
rect 41396 309134 42196 309218
rect 41396 308898 41518 309134
rect 41754 308898 41838 309134
rect 42074 308898 42196 309134
rect 41396 308866 42196 308898
rect 197872 309454 198220 309486
rect 197872 309218 197928 309454
rect 198164 309218 198220 309454
rect 197872 309134 198220 309218
rect 197872 308898 197928 309134
rect 198164 308898 198220 309134
rect 197872 308866 198220 308898
rect 292936 309454 293284 309486
rect 292936 309218 292992 309454
rect 293228 309218 293284 309454
rect 292936 309134 293284 309218
rect 292936 308898 292992 309134
rect 293228 308898 293284 309134
rect 292936 308866 293284 308898
rect 324428 309454 324776 309486
rect 324428 309218 324484 309454
rect 324720 309218 324776 309454
rect 324428 309134 324776 309218
rect 324428 308898 324484 309134
rect 324720 308898 324776 309134
rect 324428 308866 324776 308898
rect 419492 309454 419840 309486
rect 419492 309218 419548 309454
rect 419784 309218 419840 309454
rect 419492 309134 419840 309218
rect 419492 308898 419548 309134
rect 419784 308898 419840 309134
rect 419492 308866 419840 308898
rect 423100 309454 423900 309486
rect 423100 309218 423222 309454
rect 423458 309218 423542 309454
rect 423778 309218 423900 309454
rect 423100 309134 423900 309218
rect 423100 308898 423222 309134
rect 423458 308898 423542 309134
rect 423778 308898 423900 309134
rect 423100 308866 423900 308898
rect 42556 291454 43356 291486
rect 42556 291218 42678 291454
rect 42914 291218 42998 291454
rect 43234 291218 43356 291454
rect 42556 291134 43356 291218
rect 42556 290898 42678 291134
rect 42914 290898 42998 291134
rect 43234 290898 43356 291134
rect 42556 290866 43356 290898
rect 198552 291454 198900 291486
rect 198552 291218 198608 291454
rect 198844 291218 198900 291454
rect 198552 291134 198900 291218
rect 198552 290898 198608 291134
rect 198844 290898 198900 291134
rect 198552 290866 198900 290898
rect 292256 291454 292604 291486
rect 292256 291218 292312 291454
rect 292548 291218 292604 291454
rect 292256 291134 292604 291218
rect 292256 290898 292312 291134
rect 292548 290898 292604 291134
rect 292256 290866 292604 290898
rect 325108 291454 325456 291486
rect 325108 291218 325164 291454
rect 325400 291218 325456 291454
rect 325108 291134 325456 291218
rect 325108 290898 325164 291134
rect 325400 290898 325456 291134
rect 325108 290866 325456 290898
rect 418812 291454 419160 291486
rect 418812 291218 418868 291454
rect 419104 291218 419160 291454
rect 418812 291134 419160 291218
rect 418812 290898 418868 291134
rect 419104 290898 419160 291134
rect 418812 290866 419160 290898
rect 421940 291454 422740 291486
rect 421940 291218 422062 291454
rect 422298 291218 422382 291454
rect 422618 291218 422740 291454
rect 421940 291134 422740 291218
rect 421940 290898 422062 291134
rect 422298 290898 422382 291134
rect 422618 290898 422740 291134
rect 421940 290866 422740 290898
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 41396 273454 42196 273486
rect 41396 273218 41518 273454
rect 41754 273218 41838 273454
rect 42074 273218 42196 273454
rect 41396 273134 42196 273218
rect 41396 272898 41518 273134
rect 41754 272898 41838 273134
rect 42074 272898 42196 273134
rect 41396 272866 42196 272898
rect 197872 273454 198220 273486
rect 197872 273218 197928 273454
rect 198164 273218 198220 273454
rect 197872 273134 198220 273218
rect 197872 272898 197928 273134
rect 198164 272898 198220 273134
rect 197872 272866 198220 272898
rect 292936 273454 293284 273486
rect 292936 273218 292992 273454
rect 293228 273218 293284 273454
rect 292936 273134 293284 273218
rect 292936 272898 292992 273134
rect 293228 272898 293284 273134
rect 292936 272866 293284 272898
rect 324428 273454 324776 273486
rect 324428 273218 324484 273454
rect 324720 273218 324776 273454
rect 324428 273134 324776 273218
rect 324428 272898 324484 273134
rect 324720 272898 324776 273134
rect 324428 272866 324776 272898
rect 419492 273454 419840 273486
rect 419492 273218 419548 273454
rect 419784 273218 419840 273454
rect 419492 273134 419840 273218
rect 419492 272898 419548 273134
rect 419784 272898 419840 273134
rect 419492 272866 419840 272898
rect 423100 273454 423900 273486
rect 423100 273218 423222 273454
rect 423458 273218 423542 273454
rect 423778 273218 423900 273454
rect 423100 273134 423900 273218
rect 423100 272898 423222 273134
rect 423458 272898 423542 273134
rect 423778 272898 423900 273134
rect 423100 272866 423900 272898
rect 42556 255454 43356 255486
rect 42556 255218 42678 255454
rect 42914 255218 42998 255454
rect 43234 255218 43356 255454
rect 42556 255134 43356 255218
rect 42556 254898 42678 255134
rect 42914 254898 42998 255134
rect 43234 254898 43356 255134
rect 42556 254866 43356 254898
rect 421940 255454 422740 255486
rect 421940 255218 422062 255454
rect 422298 255218 422382 255454
rect 422618 255218 422740 255454
rect 421940 255134 422740 255218
rect 421940 254898 422062 255134
rect 422298 254898 422382 255134
rect 422618 254898 422740 255134
rect 421940 254866 422740 254898
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 41396 237454 42196 237486
rect 41396 237218 41518 237454
rect 41754 237218 41838 237454
rect 42074 237218 42196 237454
rect 41396 237134 42196 237218
rect 41396 236898 41518 237134
rect 41754 236898 41838 237134
rect 42074 236898 42196 237134
rect 41396 236866 42196 236898
rect 197872 237454 198220 237486
rect 197872 237218 197928 237454
rect 198164 237218 198220 237454
rect 197872 237134 198220 237218
rect 197872 236898 197928 237134
rect 198164 236898 198220 237134
rect 197872 236866 198220 236898
rect 292936 237454 293284 237486
rect 292936 237218 292992 237454
rect 293228 237218 293284 237454
rect 292936 237134 293284 237218
rect 292936 236898 292992 237134
rect 293228 236898 293284 237134
rect 292936 236866 293284 236898
rect 324428 237454 324776 237486
rect 324428 237218 324484 237454
rect 324720 237218 324776 237454
rect 324428 237134 324776 237218
rect 324428 236898 324484 237134
rect 324720 236898 324776 237134
rect 324428 236866 324776 236898
rect 419492 237454 419840 237486
rect 419492 237218 419548 237454
rect 419784 237218 419840 237454
rect 419492 237134 419840 237218
rect 419492 236898 419548 237134
rect 419784 236898 419840 237134
rect 419492 236866 419840 236898
rect 423100 237454 423900 237486
rect 423100 237218 423222 237454
rect 423458 237218 423542 237454
rect 423778 237218 423900 237454
rect 423100 237134 423900 237218
rect 423100 236898 423222 237134
rect 423458 236898 423542 237134
rect 423778 236898 423900 237134
rect 423100 236866 423900 236898
rect 42556 219454 43356 219486
rect 42556 219218 42678 219454
rect 42914 219218 42998 219454
rect 43234 219218 43356 219454
rect 42556 219134 43356 219218
rect 42556 218898 42678 219134
rect 42914 218898 42998 219134
rect 43234 218898 43356 219134
rect 42556 218866 43356 218898
rect 198552 219454 198900 219486
rect 198552 219218 198608 219454
rect 198844 219218 198900 219454
rect 198552 219134 198900 219218
rect 198552 218898 198608 219134
rect 198844 218898 198900 219134
rect 198552 218866 198900 218898
rect 292256 219454 292604 219486
rect 292256 219218 292312 219454
rect 292548 219218 292604 219454
rect 292256 219134 292604 219218
rect 292256 218898 292312 219134
rect 292548 218898 292604 219134
rect 292256 218866 292604 218898
rect 325108 219454 325456 219486
rect 325108 219218 325164 219454
rect 325400 219218 325456 219454
rect 325108 219134 325456 219218
rect 325108 218898 325164 219134
rect 325400 218898 325456 219134
rect 325108 218866 325456 218898
rect 418812 219454 419160 219486
rect 418812 219218 418868 219454
rect 419104 219218 419160 219454
rect 418812 219134 419160 219218
rect 418812 218898 418868 219134
rect 419104 218898 419160 219134
rect 418812 218866 419160 218898
rect 421940 219454 422740 219486
rect 421940 219218 422062 219454
rect 422298 219218 422382 219454
rect 422618 219218 422740 219454
rect 421940 219134 422740 219218
rect 421940 218898 422062 219134
rect 422298 218898 422382 219134
rect 422618 218898 422740 219134
rect 421940 218866 422740 218898
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 41396 201454 42196 201486
rect 41396 201218 41518 201454
rect 41754 201218 41838 201454
rect 42074 201218 42196 201454
rect 41396 201134 42196 201218
rect 41396 200898 41518 201134
rect 41754 200898 41838 201134
rect 42074 200898 42196 201134
rect 41396 200866 42196 200898
rect 197872 201454 198220 201486
rect 197872 201218 197928 201454
rect 198164 201218 198220 201454
rect 197872 201134 198220 201218
rect 197872 200898 197928 201134
rect 198164 200898 198220 201134
rect 197872 200866 198220 200898
rect 292936 201454 293284 201486
rect 292936 201218 292992 201454
rect 293228 201218 293284 201454
rect 292936 201134 293284 201218
rect 292936 200898 292992 201134
rect 293228 200898 293284 201134
rect 292936 200866 293284 200898
rect 324428 201454 324776 201486
rect 324428 201218 324484 201454
rect 324720 201218 324776 201454
rect 324428 201134 324776 201218
rect 324428 200898 324484 201134
rect 324720 200898 324776 201134
rect 324428 200866 324776 200898
rect 419492 201454 419840 201486
rect 419492 201218 419548 201454
rect 419784 201218 419840 201454
rect 419492 201134 419840 201218
rect 419492 200898 419548 201134
rect 419784 200898 419840 201134
rect 419492 200866 419840 200898
rect 423100 201454 423900 201486
rect 423100 201218 423222 201454
rect 423458 201218 423542 201454
rect 423778 201218 423900 201454
rect 423100 201134 423900 201218
rect 423100 200898 423222 201134
rect 423458 200898 423542 201134
rect 423778 200898 423900 201134
rect 423100 200866 423900 200898
rect 42556 183454 43356 183486
rect 42556 183218 42678 183454
rect 42914 183218 42998 183454
rect 43234 183218 43356 183454
rect 42556 183134 43356 183218
rect 42556 182898 42678 183134
rect 42914 182898 42998 183134
rect 43234 182898 43356 183134
rect 42556 182866 43356 182898
rect 198552 183454 198900 183486
rect 198552 183218 198608 183454
rect 198844 183218 198900 183454
rect 198552 183134 198900 183218
rect 198552 182898 198608 183134
rect 198844 182898 198900 183134
rect 198552 182866 198900 182898
rect 292256 183454 292604 183486
rect 292256 183218 292312 183454
rect 292548 183218 292604 183454
rect 292256 183134 292604 183218
rect 292256 182898 292312 183134
rect 292548 182898 292604 183134
rect 292256 182866 292604 182898
rect 325108 183454 325456 183486
rect 325108 183218 325164 183454
rect 325400 183218 325456 183454
rect 325108 183134 325456 183218
rect 325108 182898 325164 183134
rect 325400 182898 325456 183134
rect 325108 182866 325456 182898
rect 418812 183454 419160 183486
rect 418812 183218 418868 183454
rect 419104 183218 419160 183454
rect 418812 183134 419160 183218
rect 418812 182898 418868 183134
rect 419104 182898 419160 183134
rect 418812 182866 419160 182898
rect 421940 183454 422740 183486
rect 421940 183218 422062 183454
rect 422298 183218 422382 183454
rect 422618 183218 422740 183454
rect 421940 183134 422740 183218
rect 421940 182898 422062 183134
rect 422298 182898 422382 183134
rect 422618 182898 422740 183134
rect 421940 182866 422740 182898
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 41396 165454 42196 165486
rect 41396 165218 41518 165454
rect 41754 165218 41838 165454
rect 42074 165218 42196 165454
rect 41396 165134 42196 165218
rect 41396 164898 41518 165134
rect 41754 164898 41838 165134
rect 42074 164898 42196 165134
rect 41396 164866 42196 164898
rect 197872 165454 198220 165486
rect 197872 165218 197928 165454
rect 198164 165218 198220 165454
rect 197872 165134 198220 165218
rect 197872 164898 197928 165134
rect 198164 164898 198220 165134
rect 197872 164866 198220 164898
rect 292936 165454 293284 165486
rect 292936 165218 292992 165454
rect 293228 165218 293284 165454
rect 292936 165134 293284 165218
rect 292936 164898 292992 165134
rect 293228 164898 293284 165134
rect 292936 164866 293284 164898
rect 324428 165454 324776 165486
rect 324428 165218 324484 165454
rect 324720 165218 324776 165454
rect 324428 165134 324776 165218
rect 324428 164898 324484 165134
rect 324720 164898 324776 165134
rect 324428 164866 324776 164898
rect 419492 165454 419840 165486
rect 419492 165218 419548 165454
rect 419784 165218 419840 165454
rect 419492 165134 419840 165218
rect 419492 164898 419548 165134
rect 419784 164898 419840 165134
rect 419492 164866 419840 164898
rect 423100 165454 423900 165486
rect 423100 165218 423222 165454
rect 423458 165218 423542 165454
rect 423778 165218 423900 165454
rect 423100 165134 423900 165218
rect 423100 164898 423222 165134
rect 423458 164898 423542 165134
rect 423778 164898 423900 165134
rect 423100 164866 423900 164898
rect 42556 147454 43356 147486
rect 42556 147218 42678 147454
rect 42914 147218 42998 147454
rect 43234 147218 43356 147454
rect 42556 147134 43356 147218
rect 42556 146898 42678 147134
rect 42914 146898 42998 147134
rect 43234 146898 43356 147134
rect 42556 146866 43356 146898
rect 421940 147454 422740 147486
rect 421940 147218 422062 147454
rect 422298 147218 422382 147454
rect 422618 147218 422740 147454
rect 421940 147134 422740 147218
rect 421940 146898 422062 147134
rect 422298 146898 422382 147134
rect 422618 146898 422740 147134
rect 421940 146866 422740 146898
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 41396 129454 42196 129486
rect 41396 129218 41518 129454
rect 41754 129218 41838 129454
rect 42074 129218 42196 129454
rect 41396 129134 42196 129218
rect 41396 128898 41518 129134
rect 41754 128898 41838 129134
rect 42074 128898 42196 129134
rect 41396 128866 42196 128898
rect 197872 129454 198220 129486
rect 197872 129218 197928 129454
rect 198164 129218 198220 129454
rect 197872 129134 198220 129218
rect 197872 128898 197928 129134
rect 198164 128898 198220 129134
rect 197872 128866 198220 128898
rect 292936 129454 293284 129486
rect 292936 129218 292992 129454
rect 293228 129218 293284 129454
rect 292936 129134 293284 129218
rect 292936 128898 292992 129134
rect 293228 128898 293284 129134
rect 292936 128866 293284 128898
rect 324428 129454 324776 129486
rect 324428 129218 324484 129454
rect 324720 129218 324776 129454
rect 324428 129134 324776 129218
rect 324428 128898 324484 129134
rect 324720 128898 324776 129134
rect 324428 128866 324776 128898
rect 419492 129454 419840 129486
rect 419492 129218 419548 129454
rect 419784 129218 419840 129454
rect 419492 129134 419840 129218
rect 419492 128898 419548 129134
rect 419784 128898 419840 129134
rect 419492 128866 419840 128898
rect 423100 129454 423900 129486
rect 423100 129218 423222 129454
rect 423458 129218 423542 129454
rect 423778 129218 423900 129454
rect 423100 129134 423900 129218
rect 423100 128898 423222 129134
rect 423458 128898 423542 129134
rect 423778 128898 423900 129134
rect 423100 128866 423900 128898
rect 42556 111454 43356 111486
rect 42556 111218 42678 111454
rect 42914 111218 42998 111454
rect 43234 111218 43356 111454
rect 42556 111134 43356 111218
rect 42556 110898 42678 111134
rect 42914 110898 42998 111134
rect 43234 110898 43356 111134
rect 42556 110866 43356 110898
rect 198552 111454 198900 111486
rect 198552 111218 198608 111454
rect 198844 111218 198900 111454
rect 198552 111134 198900 111218
rect 198552 110898 198608 111134
rect 198844 110898 198900 111134
rect 198552 110866 198900 110898
rect 292256 111454 292604 111486
rect 292256 111218 292312 111454
rect 292548 111218 292604 111454
rect 292256 111134 292604 111218
rect 292256 110898 292312 111134
rect 292548 110898 292604 111134
rect 292256 110866 292604 110898
rect 325108 111454 325456 111486
rect 325108 111218 325164 111454
rect 325400 111218 325456 111454
rect 325108 111134 325456 111218
rect 325108 110898 325164 111134
rect 325400 110898 325456 111134
rect 325108 110866 325456 110898
rect 418812 111454 419160 111486
rect 418812 111218 418868 111454
rect 419104 111218 419160 111454
rect 418812 111134 419160 111218
rect 418812 110898 418868 111134
rect 419104 110898 419160 111134
rect 418812 110866 419160 110898
rect 421940 111454 422740 111486
rect 421940 111218 422062 111454
rect 422298 111218 422382 111454
rect 422618 111218 422740 111454
rect 421940 111134 422740 111218
rect 421940 110898 422062 111134
rect 422298 110898 422382 111134
rect 422618 110898 422740 111134
rect 421940 110866 422740 110898
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 41396 93454 42196 93486
rect 41396 93218 41518 93454
rect 41754 93218 41838 93454
rect 42074 93218 42196 93454
rect 41396 93134 42196 93218
rect 41396 92898 41518 93134
rect 41754 92898 41838 93134
rect 42074 92898 42196 93134
rect 41396 92866 42196 92898
rect 197872 93454 198220 93486
rect 197872 93218 197928 93454
rect 198164 93218 198220 93454
rect 197872 93134 198220 93218
rect 197872 92898 197928 93134
rect 198164 92898 198220 93134
rect 197872 92866 198220 92898
rect 292936 93454 293284 93486
rect 292936 93218 292992 93454
rect 293228 93218 293284 93454
rect 292936 93134 293284 93218
rect 292936 92898 292992 93134
rect 293228 92898 293284 93134
rect 292936 92866 293284 92898
rect 324428 93454 324776 93486
rect 324428 93218 324484 93454
rect 324720 93218 324776 93454
rect 324428 93134 324776 93218
rect 324428 92898 324484 93134
rect 324720 92898 324776 93134
rect 324428 92866 324776 92898
rect 419492 93454 419840 93486
rect 419492 93218 419548 93454
rect 419784 93218 419840 93454
rect 419492 93134 419840 93218
rect 419492 92898 419548 93134
rect 419784 92898 419840 93134
rect 419492 92866 419840 92898
rect 423100 93454 423900 93486
rect 423100 93218 423222 93454
rect 423458 93218 423542 93454
rect 423778 93218 423900 93454
rect 423100 93134 423900 93218
rect 423100 92898 423222 93134
rect 423458 92898 423542 93134
rect 423778 92898 423900 93134
rect 423100 92866 423900 92898
rect 42556 75454 43356 75486
rect 42556 75218 42678 75454
rect 42914 75218 42998 75454
rect 43234 75218 43356 75454
rect 42556 75134 43356 75218
rect 42556 74898 42678 75134
rect 42914 74898 42998 75134
rect 43234 74898 43356 75134
rect 42556 74866 43356 74898
rect 198552 75454 198900 75486
rect 198552 75218 198608 75454
rect 198844 75218 198900 75454
rect 198552 75134 198900 75218
rect 198552 74898 198608 75134
rect 198844 74898 198900 75134
rect 198552 74866 198900 74898
rect 292256 75454 292604 75486
rect 292256 75218 292312 75454
rect 292548 75218 292604 75454
rect 292256 75134 292604 75218
rect 292256 74898 292312 75134
rect 292548 74898 292604 75134
rect 292256 74866 292604 74898
rect 325108 75454 325456 75486
rect 325108 75218 325164 75454
rect 325400 75218 325456 75454
rect 325108 75134 325456 75218
rect 325108 74898 325164 75134
rect 325400 74898 325456 75134
rect 325108 74866 325456 74898
rect 418812 75454 419160 75486
rect 418812 75218 418868 75454
rect 419104 75218 419160 75454
rect 418812 75134 419160 75218
rect 418812 74898 418868 75134
rect 419104 74898 419160 75134
rect 418812 74866 419160 74898
rect 421940 75454 422740 75486
rect 421940 75218 422062 75454
rect 422298 75218 422382 75454
rect 422618 75218 422740 75454
rect 421940 75134 422740 75218
rect 421940 74898 422062 75134
rect 422298 74898 422382 75134
rect 422618 74898 422740 75134
rect 421940 74866 422740 74898
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 41396 57454 42196 57486
rect 41396 57218 41518 57454
rect 41754 57218 41838 57454
rect 42074 57218 42196 57454
rect 41396 57134 42196 57218
rect 41396 56898 41518 57134
rect 41754 56898 41838 57134
rect 42074 56898 42196 57134
rect 41396 56866 42196 56898
rect 197872 57454 198220 57486
rect 197872 57218 197928 57454
rect 198164 57218 198220 57454
rect 197872 57134 198220 57218
rect 197872 56898 197928 57134
rect 198164 56898 198220 57134
rect 197872 56866 198220 56898
rect 292936 57454 293284 57486
rect 292936 57218 292992 57454
rect 293228 57218 293284 57454
rect 292936 57134 293284 57218
rect 292936 56898 292992 57134
rect 293228 56898 293284 57134
rect 292936 56866 293284 56898
rect 324428 57454 324776 57486
rect 324428 57218 324484 57454
rect 324720 57218 324776 57454
rect 324428 57134 324776 57218
rect 324428 56898 324484 57134
rect 324720 56898 324776 57134
rect 324428 56866 324776 56898
rect 419492 57454 419840 57486
rect 419492 57218 419548 57454
rect 419784 57218 419840 57454
rect 419492 57134 419840 57218
rect 419492 56898 419548 57134
rect 419784 56898 419840 57134
rect 419492 56866 419840 56898
rect 423100 57454 423900 57486
rect 423100 57218 423222 57454
rect 423458 57218 423542 57454
rect 423778 57218 423900 57454
rect 423100 57134 423900 57218
rect 423100 56898 423222 57134
rect 423458 56898 423542 57134
rect 423778 56898 423900 57134
rect 423100 56866 423900 56898
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 3454 38414 38000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 38000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 38000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 38000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 38000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 38000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 38000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 38000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 3454 74414 38000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 38000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 38000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 38000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 38000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 38000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 38000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 38000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 3454 110414 38000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 38000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 38000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 38000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 38000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 38000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 38000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 38000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 3454 146414 38000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 38000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 38000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 38000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 38000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 38000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 38000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 38000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 3454 182414 38000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 38000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 38000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 38000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 38000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 38000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 38000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 38000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 3454 218414 38000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 38000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 38000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 38000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 38000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 38000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 38000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 38000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 3454 254414 38000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 38000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 38000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 38000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 38000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 38000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 38000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 38000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 3454 290414 38000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 38000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 38000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 38000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 38000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 38000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 38000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 38000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 3454 326414 38000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 38000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 38000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 38000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 38000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 38000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 38000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 38000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 3454 362414 38000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 38000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 38000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 38000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 38000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 38000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 38000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 38000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 3454 398414 38000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 38000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 38000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 38000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 38000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 38000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 38000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 38000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 42678 543218 42914 543454
rect 42998 543218 43234 543454
rect 42678 542898 42914 543134
rect 42998 542898 43234 543134
rect 200609 543218 200845 543454
rect 200609 542898 200845 543134
rect 416997 543218 417233 543454
rect 416997 542898 417233 543134
rect 422062 543218 422298 543454
rect 422382 543218 422618 543454
rect 422062 542898 422298 543134
rect 422382 542898 422618 543134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 41518 525218 41754 525454
rect 41838 525218 42074 525454
rect 41518 524898 41754 525134
rect 41838 524898 42074 525134
rect 199849 525218 200085 525454
rect 199849 524898 200085 525134
rect 205037 525218 205273 525454
rect 205037 524898 205273 525134
rect 300101 525218 300337 525454
rect 300101 524898 300337 525134
rect 317465 525218 317701 525454
rect 317465 524898 317701 525134
rect 412529 525218 412765 525454
rect 412529 524898 412765 525134
rect 417757 525218 417993 525454
rect 417757 524898 417993 525134
rect 423222 525218 423458 525454
rect 423542 525218 423778 525454
rect 423222 524898 423458 525134
rect 423542 524898 423778 525134
rect 42678 507218 42914 507454
rect 42998 507218 43234 507454
rect 42678 506898 42914 507134
rect 42998 506898 43234 507134
rect 200609 507218 200845 507454
rect 200609 506898 200845 507134
rect 205717 507218 205953 507454
rect 205717 506898 205953 507134
rect 299421 507218 299657 507454
rect 299421 506898 299657 507134
rect 318145 507218 318381 507454
rect 318145 506898 318381 507134
rect 411849 507218 412085 507454
rect 411849 506898 412085 507134
rect 416997 507218 417233 507454
rect 416997 506898 417233 507134
rect 422062 507218 422298 507454
rect 422382 507218 422618 507454
rect 422062 506898 422298 507134
rect 422382 506898 422618 507134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 41518 489218 41754 489454
rect 41838 489218 42074 489454
rect 41518 488898 41754 489134
rect 41838 488898 42074 489134
rect 199849 489218 200085 489454
rect 199849 488898 200085 489134
rect 205037 489218 205273 489454
rect 205037 488898 205273 489134
rect 300101 489218 300337 489454
rect 300101 488898 300337 489134
rect 317465 489218 317701 489454
rect 317465 488898 317701 489134
rect 412529 489218 412765 489454
rect 412529 488898 412765 489134
rect 417757 489218 417993 489454
rect 417757 488898 417993 489134
rect 423222 489218 423458 489454
rect 423542 489218 423778 489454
rect 423222 488898 423458 489134
rect 423542 488898 423778 489134
rect 42678 471218 42914 471454
rect 42998 471218 43234 471454
rect 42678 470898 42914 471134
rect 42998 470898 43234 471134
rect 200609 471218 200845 471454
rect 200609 470898 200845 471134
rect 205717 471218 205953 471454
rect 205717 470898 205953 471134
rect 299421 471218 299657 471454
rect 299421 470898 299657 471134
rect 318145 471218 318381 471454
rect 318145 470898 318381 471134
rect 411849 471218 412085 471454
rect 411849 470898 412085 471134
rect 416997 471218 417233 471454
rect 416997 470898 417233 471134
rect 422062 471218 422298 471454
rect 422382 471218 422618 471454
rect 422062 470898 422298 471134
rect 422382 470898 422618 471134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 41518 453218 41754 453454
rect 41838 453218 42074 453454
rect 41518 452898 41754 453134
rect 41838 452898 42074 453134
rect 423222 453218 423458 453454
rect 423542 453218 423778 453454
rect 423222 452898 423458 453134
rect 423542 452898 423778 453134
rect 42678 435218 42914 435454
rect 42998 435218 43234 435454
rect 42678 434898 42914 435134
rect 42998 434898 43234 435134
rect 198608 435218 198844 435454
rect 198608 434898 198844 435134
rect 292312 435218 292548 435454
rect 292312 434898 292548 435134
rect 325164 435218 325400 435454
rect 325164 434898 325400 435134
rect 418868 435218 419104 435454
rect 418868 434898 419104 435134
rect 422062 435218 422298 435454
rect 422382 435218 422618 435454
rect 422062 434898 422298 435134
rect 422382 434898 422618 435134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 41518 417218 41754 417454
rect 41838 417218 42074 417454
rect 41518 416898 41754 417134
rect 41838 416898 42074 417134
rect 197928 417218 198164 417454
rect 197928 416898 198164 417134
rect 292992 417218 293228 417454
rect 292992 416898 293228 417134
rect 324484 417218 324720 417454
rect 324484 416898 324720 417134
rect 419548 417218 419784 417454
rect 419548 416898 419784 417134
rect 423222 417218 423458 417454
rect 423542 417218 423778 417454
rect 423222 416898 423458 417134
rect 423542 416898 423778 417134
rect 42678 399218 42914 399454
rect 42998 399218 43234 399454
rect 42678 398898 42914 399134
rect 42998 398898 43234 399134
rect 198608 399218 198844 399454
rect 198608 398898 198844 399134
rect 292312 399218 292548 399454
rect 292312 398898 292548 399134
rect 325164 399218 325400 399454
rect 325164 398898 325400 399134
rect 418868 399218 419104 399454
rect 418868 398898 419104 399134
rect 422062 399218 422298 399454
rect 422382 399218 422618 399454
rect 422062 398898 422298 399134
rect 422382 398898 422618 399134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 41518 381218 41754 381454
rect 41838 381218 42074 381454
rect 41518 380898 41754 381134
rect 41838 380898 42074 381134
rect 197928 381218 198164 381454
rect 197928 380898 198164 381134
rect 292992 381218 293228 381454
rect 292992 380898 293228 381134
rect 324484 381218 324720 381454
rect 324484 380898 324720 381134
rect 419548 381218 419784 381454
rect 419548 380898 419784 381134
rect 423222 381218 423458 381454
rect 423542 381218 423778 381454
rect 423222 380898 423458 381134
rect 423542 380898 423778 381134
rect 42678 363218 42914 363454
rect 42998 363218 43234 363454
rect 42678 362898 42914 363134
rect 42998 362898 43234 363134
rect 422062 363218 422298 363454
rect 422382 363218 422618 363454
rect 422062 362898 422298 363134
rect 422382 362898 422618 363134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 41518 345218 41754 345454
rect 41838 345218 42074 345454
rect 41518 344898 41754 345134
rect 41838 344898 42074 345134
rect 423222 345218 423458 345454
rect 423542 345218 423778 345454
rect 423222 344898 423458 345134
rect 423542 344898 423778 345134
rect 42678 327218 42914 327454
rect 42998 327218 43234 327454
rect 42678 326898 42914 327134
rect 42998 326898 43234 327134
rect 198608 327218 198844 327454
rect 198608 326898 198844 327134
rect 292312 327218 292548 327454
rect 292312 326898 292548 327134
rect 325164 327218 325400 327454
rect 325164 326898 325400 327134
rect 418868 327218 419104 327454
rect 418868 326898 419104 327134
rect 422062 327218 422298 327454
rect 422382 327218 422618 327454
rect 422062 326898 422298 327134
rect 422382 326898 422618 327134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 41518 309218 41754 309454
rect 41838 309218 42074 309454
rect 41518 308898 41754 309134
rect 41838 308898 42074 309134
rect 197928 309218 198164 309454
rect 197928 308898 198164 309134
rect 292992 309218 293228 309454
rect 292992 308898 293228 309134
rect 324484 309218 324720 309454
rect 324484 308898 324720 309134
rect 419548 309218 419784 309454
rect 419548 308898 419784 309134
rect 423222 309218 423458 309454
rect 423542 309218 423778 309454
rect 423222 308898 423458 309134
rect 423542 308898 423778 309134
rect 42678 291218 42914 291454
rect 42998 291218 43234 291454
rect 42678 290898 42914 291134
rect 42998 290898 43234 291134
rect 198608 291218 198844 291454
rect 198608 290898 198844 291134
rect 292312 291218 292548 291454
rect 292312 290898 292548 291134
rect 325164 291218 325400 291454
rect 325164 290898 325400 291134
rect 418868 291218 419104 291454
rect 418868 290898 419104 291134
rect 422062 291218 422298 291454
rect 422382 291218 422618 291454
rect 422062 290898 422298 291134
rect 422382 290898 422618 291134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 41518 273218 41754 273454
rect 41838 273218 42074 273454
rect 41518 272898 41754 273134
rect 41838 272898 42074 273134
rect 197928 273218 198164 273454
rect 197928 272898 198164 273134
rect 292992 273218 293228 273454
rect 292992 272898 293228 273134
rect 324484 273218 324720 273454
rect 324484 272898 324720 273134
rect 419548 273218 419784 273454
rect 419548 272898 419784 273134
rect 423222 273218 423458 273454
rect 423542 273218 423778 273454
rect 423222 272898 423458 273134
rect 423542 272898 423778 273134
rect 42678 255218 42914 255454
rect 42998 255218 43234 255454
rect 42678 254898 42914 255134
rect 42998 254898 43234 255134
rect 422062 255218 422298 255454
rect 422382 255218 422618 255454
rect 422062 254898 422298 255134
rect 422382 254898 422618 255134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 41518 237218 41754 237454
rect 41838 237218 42074 237454
rect 41518 236898 41754 237134
rect 41838 236898 42074 237134
rect 197928 237218 198164 237454
rect 197928 236898 198164 237134
rect 292992 237218 293228 237454
rect 292992 236898 293228 237134
rect 324484 237218 324720 237454
rect 324484 236898 324720 237134
rect 419548 237218 419784 237454
rect 419548 236898 419784 237134
rect 423222 237218 423458 237454
rect 423542 237218 423778 237454
rect 423222 236898 423458 237134
rect 423542 236898 423778 237134
rect 42678 219218 42914 219454
rect 42998 219218 43234 219454
rect 42678 218898 42914 219134
rect 42998 218898 43234 219134
rect 198608 219218 198844 219454
rect 198608 218898 198844 219134
rect 292312 219218 292548 219454
rect 292312 218898 292548 219134
rect 325164 219218 325400 219454
rect 325164 218898 325400 219134
rect 418868 219218 419104 219454
rect 418868 218898 419104 219134
rect 422062 219218 422298 219454
rect 422382 219218 422618 219454
rect 422062 218898 422298 219134
rect 422382 218898 422618 219134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 41518 201218 41754 201454
rect 41838 201218 42074 201454
rect 41518 200898 41754 201134
rect 41838 200898 42074 201134
rect 197928 201218 198164 201454
rect 197928 200898 198164 201134
rect 292992 201218 293228 201454
rect 292992 200898 293228 201134
rect 324484 201218 324720 201454
rect 324484 200898 324720 201134
rect 419548 201218 419784 201454
rect 419548 200898 419784 201134
rect 423222 201218 423458 201454
rect 423542 201218 423778 201454
rect 423222 200898 423458 201134
rect 423542 200898 423778 201134
rect 42678 183218 42914 183454
rect 42998 183218 43234 183454
rect 42678 182898 42914 183134
rect 42998 182898 43234 183134
rect 198608 183218 198844 183454
rect 198608 182898 198844 183134
rect 292312 183218 292548 183454
rect 292312 182898 292548 183134
rect 325164 183218 325400 183454
rect 325164 182898 325400 183134
rect 418868 183218 419104 183454
rect 418868 182898 419104 183134
rect 422062 183218 422298 183454
rect 422382 183218 422618 183454
rect 422062 182898 422298 183134
rect 422382 182898 422618 183134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 41518 165218 41754 165454
rect 41838 165218 42074 165454
rect 41518 164898 41754 165134
rect 41838 164898 42074 165134
rect 197928 165218 198164 165454
rect 197928 164898 198164 165134
rect 292992 165218 293228 165454
rect 292992 164898 293228 165134
rect 324484 165218 324720 165454
rect 324484 164898 324720 165134
rect 419548 165218 419784 165454
rect 419548 164898 419784 165134
rect 423222 165218 423458 165454
rect 423542 165218 423778 165454
rect 423222 164898 423458 165134
rect 423542 164898 423778 165134
rect 42678 147218 42914 147454
rect 42998 147218 43234 147454
rect 42678 146898 42914 147134
rect 42998 146898 43234 147134
rect 422062 147218 422298 147454
rect 422382 147218 422618 147454
rect 422062 146898 422298 147134
rect 422382 146898 422618 147134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 41518 129218 41754 129454
rect 41838 129218 42074 129454
rect 41518 128898 41754 129134
rect 41838 128898 42074 129134
rect 197928 129218 198164 129454
rect 197928 128898 198164 129134
rect 292992 129218 293228 129454
rect 292992 128898 293228 129134
rect 324484 129218 324720 129454
rect 324484 128898 324720 129134
rect 419548 129218 419784 129454
rect 419548 128898 419784 129134
rect 423222 129218 423458 129454
rect 423542 129218 423778 129454
rect 423222 128898 423458 129134
rect 423542 128898 423778 129134
rect 42678 111218 42914 111454
rect 42998 111218 43234 111454
rect 42678 110898 42914 111134
rect 42998 110898 43234 111134
rect 198608 111218 198844 111454
rect 198608 110898 198844 111134
rect 292312 111218 292548 111454
rect 292312 110898 292548 111134
rect 325164 111218 325400 111454
rect 325164 110898 325400 111134
rect 418868 111218 419104 111454
rect 418868 110898 419104 111134
rect 422062 111218 422298 111454
rect 422382 111218 422618 111454
rect 422062 110898 422298 111134
rect 422382 110898 422618 111134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 41518 93218 41754 93454
rect 41838 93218 42074 93454
rect 41518 92898 41754 93134
rect 41838 92898 42074 93134
rect 197928 93218 198164 93454
rect 197928 92898 198164 93134
rect 292992 93218 293228 93454
rect 292992 92898 293228 93134
rect 324484 93218 324720 93454
rect 324484 92898 324720 93134
rect 419548 93218 419784 93454
rect 419548 92898 419784 93134
rect 423222 93218 423458 93454
rect 423542 93218 423778 93454
rect 423222 92898 423458 93134
rect 423542 92898 423778 93134
rect 42678 75218 42914 75454
rect 42998 75218 43234 75454
rect 42678 74898 42914 75134
rect 42998 74898 43234 75134
rect 198608 75218 198844 75454
rect 198608 74898 198844 75134
rect 292312 75218 292548 75454
rect 292312 74898 292548 75134
rect 325164 75218 325400 75454
rect 325164 74898 325400 75134
rect 418868 75218 419104 75454
rect 418868 74898 419104 75134
rect 422062 75218 422298 75454
rect 422382 75218 422618 75454
rect 422062 74898 422298 75134
rect 422382 74898 422618 75134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 41518 57218 41754 57454
rect 41838 57218 42074 57454
rect 41518 56898 41754 57134
rect 41838 56898 42074 57134
rect 197928 57218 198164 57454
rect 197928 56898 198164 57134
rect 292992 57218 293228 57454
rect 292992 56898 293228 57134
rect 324484 57218 324720 57454
rect 324484 56898 324720 57134
rect 419548 57218 419784 57454
rect 419548 56898 419784 57134
rect 423222 57218 423458 57454
rect 423542 57218 423778 57454
rect 423222 56898 423458 57134
rect 423542 56898 423778 57134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 42678 543454
rect 42914 543218 42998 543454
rect 43234 543218 200609 543454
rect 200845 543218 416997 543454
rect 417233 543218 422062 543454
rect 422298 543218 422382 543454
rect 422618 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 42678 543134
rect 42914 542898 42998 543134
rect 43234 542898 200609 543134
rect 200845 542898 416997 543134
rect 417233 542898 422062 543134
rect 422298 542898 422382 543134
rect 422618 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 41518 525454
rect 41754 525218 41838 525454
rect 42074 525218 199849 525454
rect 200085 525218 205037 525454
rect 205273 525218 300101 525454
rect 300337 525218 317465 525454
rect 317701 525218 412529 525454
rect 412765 525218 417757 525454
rect 417993 525218 423222 525454
rect 423458 525218 423542 525454
rect 423778 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 41518 525134
rect 41754 524898 41838 525134
rect 42074 524898 199849 525134
rect 200085 524898 205037 525134
rect 205273 524898 300101 525134
rect 300337 524898 317465 525134
rect 317701 524898 412529 525134
rect 412765 524898 417757 525134
rect 417993 524898 423222 525134
rect 423458 524898 423542 525134
rect 423778 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 42678 507454
rect 42914 507218 42998 507454
rect 43234 507218 200609 507454
rect 200845 507218 205717 507454
rect 205953 507218 299421 507454
rect 299657 507218 318145 507454
rect 318381 507218 411849 507454
rect 412085 507218 416997 507454
rect 417233 507218 422062 507454
rect 422298 507218 422382 507454
rect 422618 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 42678 507134
rect 42914 506898 42998 507134
rect 43234 506898 200609 507134
rect 200845 506898 205717 507134
rect 205953 506898 299421 507134
rect 299657 506898 318145 507134
rect 318381 506898 411849 507134
rect 412085 506898 416997 507134
rect 417233 506898 422062 507134
rect 422298 506898 422382 507134
rect 422618 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 41518 489454
rect 41754 489218 41838 489454
rect 42074 489218 199849 489454
rect 200085 489218 205037 489454
rect 205273 489218 300101 489454
rect 300337 489218 317465 489454
rect 317701 489218 412529 489454
rect 412765 489218 417757 489454
rect 417993 489218 423222 489454
rect 423458 489218 423542 489454
rect 423778 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 41518 489134
rect 41754 488898 41838 489134
rect 42074 488898 199849 489134
rect 200085 488898 205037 489134
rect 205273 488898 300101 489134
rect 300337 488898 317465 489134
rect 317701 488898 412529 489134
rect 412765 488898 417757 489134
rect 417993 488898 423222 489134
rect 423458 488898 423542 489134
rect 423778 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 42678 471454
rect 42914 471218 42998 471454
rect 43234 471218 200609 471454
rect 200845 471218 205717 471454
rect 205953 471218 299421 471454
rect 299657 471218 318145 471454
rect 318381 471218 411849 471454
rect 412085 471218 416997 471454
rect 417233 471218 422062 471454
rect 422298 471218 422382 471454
rect 422618 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 42678 471134
rect 42914 470898 42998 471134
rect 43234 470898 200609 471134
rect 200845 470898 205717 471134
rect 205953 470898 299421 471134
rect 299657 470898 318145 471134
rect 318381 470898 411849 471134
rect 412085 470898 416997 471134
rect 417233 470898 422062 471134
rect 422298 470898 422382 471134
rect 422618 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 41518 453454
rect 41754 453218 41838 453454
rect 42074 453218 423222 453454
rect 423458 453218 423542 453454
rect 423778 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 41518 453134
rect 41754 452898 41838 453134
rect 42074 452898 423222 453134
rect 423458 452898 423542 453134
rect 423778 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 42678 435454
rect 42914 435218 42998 435454
rect 43234 435218 198608 435454
rect 198844 435218 292312 435454
rect 292548 435218 325164 435454
rect 325400 435218 418868 435454
rect 419104 435218 422062 435454
rect 422298 435218 422382 435454
rect 422618 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 42678 435134
rect 42914 434898 42998 435134
rect 43234 434898 198608 435134
rect 198844 434898 292312 435134
rect 292548 434898 325164 435134
rect 325400 434898 418868 435134
rect 419104 434898 422062 435134
rect 422298 434898 422382 435134
rect 422618 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 41518 417454
rect 41754 417218 41838 417454
rect 42074 417218 197928 417454
rect 198164 417218 292992 417454
rect 293228 417218 324484 417454
rect 324720 417218 419548 417454
rect 419784 417218 423222 417454
rect 423458 417218 423542 417454
rect 423778 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 41518 417134
rect 41754 416898 41838 417134
rect 42074 416898 197928 417134
rect 198164 416898 292992 417134
rect 293228 416898 324484 417134
rect 324720 416898 419548 417134
rect 419784 416898 423222 417134
rect 423458 416898 423542 417134
rect 423778 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 42678 399454
rect 42914 399218 42998 399454
rect 43234 399218 198608 399454
rect 198844 399218 292312 399454
rect 292548 399218 325164 399454
rect 325400 399218 418868 399454
rect 419104 399218 422062 399454
rect 422298 399218 422382 399454
rect 422618 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 42678 399134
rect 42914 398898 42998 399134
rect 43234 398898 198608 399134
rect 198844 398898 292312 399134
rect 292548 398898 325164 399134
rect 325400 398898 418868 399134
rect 419104 398898 422062 399134
rect 422298 398898 422382 399134
rect 422618 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 41518 381454
rect 41754 381218 41838 381454
rect 42074 381218 197928 381454
rect 198164 381218 292992 381454
rect 293228 381218 324484 381454
rect 324720 381218 419548 381454
rect 419784 381218 423222 381454
rect 423458 381218 423542 381454
rect 423778 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 41518 381134
rect 41754 380898 41838 381134
rect 42074 380898 197928 381134
rect 198164 380898 292992 381134
rect 293228 380898 324484 381134
rect 324720 380898 419548 381134
rect 419784 380898 423222 381134
rect 423458 380898 423542 381134
rect 423778 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 42678 363454
rect 42914 363218 42998 363454
rect 43234 363218 422062 363454
rect 422298 363218 422382 363454
rect 422618 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 42678 363134
rect 42914 362898 42998 363134
rect 43234 362898 422062 363134
rect 422298 362898 422382 363134
rect 422618 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 41518 345454
rect 41754 345218 41838 345454
rect 42074 345218 423222 345454
rect 423458 345218 423542 345454
rect 423778 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 41518 345134
rect 41754 344898 41838 345134
rect 42074 344898 423222 345134
rect 423458 344898 423542 345134
rect 423778 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 42678 327454
rect 42914 327218 42998 327454
rect 43234 327218 198608 327454
rect 198844 327218 292312 327454
rect 292548 327218 325164 327454
rect 325400 327218 418868 327454
rect 419104 327218 422062 327454
rect 422298 327218 422382 327454
rect 422618 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 42678 327134
rect 42914 326898 42998 327134
rect 43234 326898 198608 327134
rect 198844 326898 292312 327134
rect 292548 326898 325164 327134
rect 325400 326898 418868 327134
rect 419104 326898 422062 327134
rect 422298 326898 422382 327134
rect 422618 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 41518 309454
rect 41754 309218 41838 309454
rect 42074 309218 197928 309454
rect 198164 309218 292992 309454
rect 293228 309218 324484 309454
rect 324720 309218 419548 309454
rect 419784 309218 423222 309454
rect 423458 309218 423542 309454
rect 423778 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 41518 309134
rect 41754 308898 41838 309134
rect 42074 308898 197928 309134
rect 198164 308898 292992 309134
rect 293228 308898 324484 309134
rect 324720 308898 419548 309134
rect 419784 308898 423222 309134
rect 423458 308898 423542 309134
rect 423778 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 42678 291454
rect 42914 291218 42998 291454
rect 43234 291218 198608 291454
rect 198844 291218 292312 291454
rect 292548 291218 325164 291454
rect 325400 291218 418868 291454
rect 419104 291218 422062 291454
rect 422298 291218 422382 291454
rect 422618 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 42678 291134
rect 42914 290898 42998 291134
rect 43234 290898 198608 291134
rect 198844 290898 292312 291134
rect 292548 290898 325164 291134
rect 325400 290898 418868 291134
rect 419104 290898 422062 291134
rect 422298 290898 422382 291134
rect 422618 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 41518 273454
rect 41754 273218 41838 273454
rect 42074 273218 197928 273454
rect 198164 273218 292992 273454
rect 293228 273218 324484 273454
rect 324720 273218 419548 273454
rect 419784 273218 423222 273454
rect 423458 273218 423542 273454
rect 423778 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 41518 273134
rect 41754 272898 41838 273134
rect 42074 272898 197928 273134
rect 198164 272898 292992 273134
rect 293228 272898 324484 273134
rect 324720 272898 419548 273134
rect 419784 272898 423222 273134
rect 423458 272898 423542 273134
rect 423778 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 42678 255454
rect 42914 255218 42998 255454
rect 43234 255218 422062 255454
rect 422298 255218 422382 255454
rect 422618 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 42678 255134
rect 42914 254898 42998 255134
rect 43234 254898 422062 255134
rect 422298 254898 422382 255134
rect 422618 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 41518 237454
rect 41754 237218 41838 237454
rect 42074 237218 197928 237454
rect 198164 237218 292992 237454
rect 293228 237218 324484 237454
rect 324720 237218 419548 237454
rect 419784 237218 423222 237454
rect 423458 237218 423542 237454
rect 423778 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 41518 237134
rect 41754 236898 41838 237134
rect 42074 236898 197928 237134
rect 198164 236898 292992 237134
rect 293228 236898 324484 237134
rect 324720 236898 419548 237134
rect 419784 236898 423222 237134
rect 423458 236898 423542 237134
rect 423778 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 42678 219454
rect 42914 219218 42998 219454
rect 43234 219218 198608 219454
rect 198844 219218 292312 219454
rect 292548 219218 325164 219454
rect 325400 219218 418868 219454
rect 419104 219218 422062 219454
rect 422298 219218 422382 219454
rect 422618 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 42678 219134
rect 42914 218898 42998 219134
rect 43234 218898 198608 219134
rect 198844 218898 292312 219134
rect 292548 218898 325164 219134
rect 325400 218898 418868 219134
rect 419104 218898 422062 219134
rect 422298 218898 422382 219134
rect 422618 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 41518 201454
rect 41754 201218 41838 201454
rect 42074 201218 197928 201454
rect 198164 201218 292992 201454
rect 293228 201218 324484 201454
rect 324720 201218 419548 201454
rect 419784 201218 423222 201454
rect 423458 201218 423542 201454
rect 423778 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 41518 201134
rect 41754 200898 41838 201134
rect 42074 200898 197928 201134
rect 198164 200898 292992 201134
rect 293228 200898 324484 201134
rect 324720 200898 419548 201134
rect 419784 200898 423222 201134
rect 423458 200898 423542 201134
rect 423778 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 42678 183454
rect 42914 183218 42998 183454
rect 43234 183218 198608 183454
rect 198844 183218 292312 183454
rect 292548 183218 325164 183454
rect 325400 183218 418868 183454
rect 419104 183218 422062 183454
rect 422298 183218 422382 183454
rect 422618 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 42678 183134
rect 42914 182898 42998 183134
rect 43234 182898 198608 183134
rect 198844 182898 292312 183134
rect 292548 182898 325164 183134
rect 325400 182898 418868 183134
rect 419104 182898 422062 183134
rect 422298 182898 422382 183134
rect 422618 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 41518 165454
rect 41754 165218 41838 165454
rect 42074 165218 197928 165454
rect 198164 165218 292992 165454
rect 293228 165218 324484 165454
rect 324720 165218 419548 165454
rect 419784 165218 423222 165454
rect 423458 165218 423542 165454
rect 423778 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 41518 165134
rect 41754 164898 41838 165134
rect 42074 164898 197928 165134
rect 198164 164898 292992 165134
rect 293228 164898 324484 165134
rect 324720 164898 419548 165134
rect 419784 164898 423222 165134
rect 423458 164898 423542 165134
rect 423778 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 42678 147454
rect 42914 147218 42998 147454
rect 43234 147218 422062 147454
rect 422298 147218 422382 147454
rect 422618 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 42678 147134
rect 42914 146898 42998 147134
rect 43234 146898 422062 147134
rect 422298 146898 422382 147134
rect 422618 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 41518 129454
rect 41754 129218 41838 129454
rect 42074 129218 197928 129454
rect 198164 129218 292992 129454
rect 293228 129218 324484 129454
rect 324720 129218 419548 129454
rect 419784 129218 423222 129454
rect 423458 129218 423542 129454
rect 423778 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 41518 129134
rect 41754 128898 41838 129134
rect 42074 128898 197928 129134
rect 198164 128898 292992 129134
rect 293228 128898 324484 129134
rect 324720 128898 419548 129134
rect 419784 128898 423222 129134
rect 423458 128898 423542 129134
rect 423778 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 42678 111454
rect 42914 111218 42998 111454
rect 43234 111218 198608 111454
rect 198844 111218 292312 111454
rect 292548 111218 325164 111454
rect 325400 111218 418868 111454
rect 419104 111218 422062 111454
rect 422298 111218 422382 111454
rect 422618 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 42678 111134
rect 42914 110898 42998 111134
rect 43234 110898 198608 111134
rect 198844 110898 292312 111134
rect 292548 110898 325164 111134
rect 325400 110898 418868 111134
rect 419104 110898 422062 111134
rect 422298 110898 422382 111134
rect 422618 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 41518 93454
rect 41754 93218 41838 93454
rect 42074 93218 197928 93454
rect 198164 93218 292992 93454
rect 293228 93218 324484 93454
rect 324720 93218 419548 93454
rect 419784 93218 423222 93454
rect 423458 93218 423542 93454
rect 423778 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 41518 93134
rect 41754 92898 41838 93134
rect 42074 92898 197928 93134
rect 198164 92898 292992 93134
rect 293228 92898 324484 93134
rect 324720 92898 419548 93134
rect 419784 92898 423222 93134
rect 423458 92898 423542 93134
rect 423778 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 42678 75454
rect 42914 75218 42998 75454
rect 43234 75218 198608 75454
rect 198844 75218 292312 75454
rect 292548 75218 325164 75454
rect 325400 75218 418868 75454
rect 419104 75218 422062 75454
rect 422298 75218 422382 75454
rect 422618 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 42678 75134
rect 42914 74898 42998 75134
rect 43234 74898 198608 75134
rect 198844 74898 292312 75134
rect 292548 74898 325164 75134
rect 325400 74898 418868 75134
rect 419104 74898 422062 75134
rect 422298 74898 422382 75134
rect 422618 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 41518 57454
rect 41754 57218 41838 57454
rect 42074 57218 197928 57454
rect 198164 57218 292992 57454
rect 293228 57218 324484 57454
rect 324720 57218 419548 57454
rect 419784 57218 423222 57454
rect 423458 57218 423542 57454
rect 423778 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 41518 57134
rect 41754 56898 41838 57134
rect 42074 56898 197928 57134
rect 198164 56898 292992 57134
rect 293228 56898 324484 57134
rect 324720 56898 419548 57134
rect 419784 56898 423222 57134
rect 423458 56898 423542 57134
rect 423778 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rest_top  mprj
timestamp 0
transform 1 0 40000 0 1 40000
box 0 0 385296 519044
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 38000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 561044 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 561044 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 561044 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 561044 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 561044 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 561044 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 561044 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 561044 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 561044 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 561044 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 561044 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 38000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 561044 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 561044 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 561044 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 561044 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 561044 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 561044 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 561044 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 561044 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 561044 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 561044 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 561044 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 38000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 561044 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 561044 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 561044 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 561044 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 561044 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 561044 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 561044 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 561044 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 561044 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 561044 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 561044 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 38000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 561044 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 561044 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 561044 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 561044 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 561044 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 561044 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 561044 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 561044 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 561044 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 561044 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 561044 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 38000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 561044 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 561044 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 561044 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 561044 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 561044 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 561044 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 561044 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 561044 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 561044 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 561044 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 561044 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 38000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 561044 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 561044 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 561044 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 561044 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 561044 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 561044 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 561044 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 561044 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 561044 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 561044 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 561044 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 38000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 561044 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 561044 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 561044 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 561044 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 561044 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 561044 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 561044 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 561044 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 561044 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 561044 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 561044 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 38000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 561044 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 561044 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 561044 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 561044 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 561044 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 561044 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 561044 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 561044 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 561044 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 561044 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 561044 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
